// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/fuji/X_GTXE2_CHANNEL.v,v 1.11 2010/10/01 14:17:17 vandanad Exp $
///////////////////////////////////////////////////////
//  Copyright (c) 2010 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     : 13.0.1
//  \  \           Description : Xilinx Functional Simulation Library Component
//  /  /                      
// /__/   /\       Filename    : X_GTXE2_CHANNEL.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Revision:		1.0
//  11/10/09 - CR - Initial version
//  11/20/09 - CR - Attribute updates in YML
//  04/27/10 - CR - YML update
//  05/26/10 - CR561562 - SATA_CPLL_CFG attribute bug fixed
//  06/10/10 - CR564909 - publish complete verilog unisim wrapper
//  06/17/10 - CR564909 - YML & RTL updates
//  06/17/10 - CR564909 - YML & RTL updates
//  08/05/10 - CR569019 - GTXE2 YML and secureip update
//  09/15/10 - CR575512 - GTXE2 YML and secureip update
/////////////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module X_GTXE2_CHANNEL (
  CPLLFBCLKLOST,
  CPLLLOCK,
  CPLLREFCLKLOST,
  DMONITOROUT,
  DRPDO,
  DRPRDY,
  EYESCANDATAERROR,
  GTREFCLKMONITOR,
  GTXTXN,
  GTXTXP,
  PCSRSVDOUT,
  PHYSTATUS,
  RXBUFSTATUS,
  RXBYTEISALIGNED,
  RXBYTEREALIGN,
  RXCDRLOCK,
  RXCHANBONDSEQ,
  RXCHANISALIGNED,
  RXCHANREALIGN,
  RXCHARISCOMMA,
  RXCHARISK,
  RXCHBONDO,
  RXCLKCORCNT,
  RXCOMINITDET,
  RXCOMMADET,
  RXCOMSASDET,
  RXCOMWAKEDET,
  RXDATA,
  RXDATAVALID,
  RXDISPERR,
  RXDLYSRESETDONE,
  RXELECIDLE,
  RXHEADER,
  RXHEADERVALID,
  RXMONITOROUT,
  RXNOTINTABLE,
  RXOUTCLK,
  RXOUTCLKFABRIC,
  RXOUTCLKPCS,
  RXPHALIGNDONE,
  RXPHMONITOR,
  RXPHSLIPMONITOR,
  RXPRBSERR,
  RXQPISENN,
  RXQPISENP,
  RXRATEDONE,
  RXRESETDONE,
  RXSTARTOFSEQ,
  RXSTATUS,
  RXVALID,
  TSTOUT,
  TXBUFSTATUS,
  TXCOMFINISH,
  TXDLYSRESETDONE,
  TXGEARBOXREADY,
  TXOUTCLK,
  TXOUTCLKFABRIC,
  TXOUTCLKPCS,
  TXPHALIGNDONE,
  TXPHINITDONE,
  TXQPISENN,
  TXQPISENP,
  TXRATEDONE,
  TXRESETDONE,

  CFGRESET,
  CLKRSVD,
  CPLLLOCKDETCLK,
  CPLLLOCKEN,
  CPLLPD,
  CPLLREFCLKSEL,
  CPLLRESET,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  EYESCANMODE,
  EYESCANRESET,
  EYESCANTRIGGER,
  GTGREFCLK,
  GTNORTHREFCLK0,
  GTNORTHREFCLK1,
  GTREFCLK0,
  GTREFCLK1,
  GTRESETSEL,
  GTRSVD,
  GTRXRESET,
  GTSOUTHREFCLK0,
  GTSOUTHREFCLK1,
  GTTXRESET,
  GTXRXN,
  GTXRXP,
  LOOPBACK,
  PCSRSVDIN,
  PCSRSVDIN2,
  PMARSVDIN,
  PMARSVDIN2,
  QPLLCLK,
  QPLLREFCLK,
  RESETOVRD,
  RX8B10BEN,
  RXBUFRESET,
  RXCDRFREQRESET,
  RXCDRHOLD,
  RXCDROVRDEN,
  RXCDRRESET,
  RXCDRRESETRSV,
  RXCHBONDEN,
  RXCHBONDI,
  RXCHBONDLEVEL,
  RXCHBONDMASTER,
  RXCHBONDSLAVE,
  RXCOMMADETEN,
  RXDDIEN,
  RXDFEAGCHOLD,
  RXDFEAGCOVRDEN,
  RXDFECM1EN,
  RXDFELFHOLD,
  RXDFELFOVRDEN,
  RXDFELPMRESET,
  RXDFETAP2HOLD,
  RXDFETAP2OVRDEN,
  RXDFETAP3HOLD,
  RXDFETAP3OVRDEN,
  RXDFETAP4HOLD,
  RXDFETAP4OVRDEN,
  RXDFETAP5HOLD,
  RXDFETAP5OVRDEN,
  RXDFEUTHOLD,
  RXDFEUTOVRDEN,
  RXDFEVPHOLD,
  RXDFEVPOVRDEN,
  RXDFEVSEN,
  RXDFEXYDEN,
  RXDFEXYDHOLD,
  RXDFEXYDOVRDEN,
  RXDLYBYPASS,
  RXDLYEN,
  RXDLYOVRDEN,
  RXDLYSRESET,
  RXELECIDLEMODE,
  RXGEARBOXSLIP,
  RXLPMEN,
  RXLPMHFHOLD,
  RXLPMHFOVRDEN,
  RXLPMLFHOLD,
  RXLPMLFKLOVRDEN,
  RXMCOMMAALIGNEN,
  RXMONITORSEL,
  RXOOBRESET,
  RXOSHOLD,
  RXOSOVRDEN,
  RXOUTCLKSEL,
  RXPCOMMAALIGNEN,
  RXPCSRESET,
  RXPD,
  RXPHALIGN,
  RXPHALIGNEN,
  RXPHDLYPD,
  RXPHDLYRESET,
  RXPHOVRDEN,
  RXPMARESET,
  RXPOLARITY,
  RXPRBSCNTRESET,
  RXPRBSSEL,
  RXQPIEN,
  RXRATE,
  RXSLIDE,
  RXSYSCLKSEL,
  RXUSERRDY,
  RXUSRCLK,
  RXUSRCLK2,
  SETERRSTATUS,
  TSTIN,
  TX8B10BBYPASS,
  TX8B10BEN,
  TXBUFDIFFCTRL,
  TXCHARDISPMODE,
  TXCHARDISPVAL,
  TXCHARISK,
  TXCOMINIT,
  TXCOMSAS,
  TXCOMWAKE,
  TXDATA,
  TXDEEMPH,
  TXDETECTRX,
  TXDIFFCTRL,
  TXDIFFPD,
  TXDLYBYPASS,
  TXDLYEN,
  TXDLYHOLD,
  TXDLYOVRDEN,
  TXDLYSRESET,
  TXDLYUPDOWN,
  TXELECIDLE,
  TXHEADER,
  TXINHIBIT,
  TXMAINCURSOR,
  TXMARGIN,
  TXOUTCLKSEL,
  TXPCSRESET,
  TXPD,
  TXPDELECIDLEMODE,
  TXPHALIGN,
  TXPHALIGNEN,
  TXPHDLYPD,
  TXPHDLYRESET,
  TXPHDLYTSTCLK,
  TXPHINIT,
  TXPHOVRDEN,
  TXPISOPD,
  TXPMARESET,
  TXPOLARITY,
  TXPOSTCURSOR,
  TXPOSTCURSORINV,
  TXPRBSFORCEERR,
  TXPRBSSEL,
  TXPRECURSOR,
  TXPRECURSORINV,
  TXQPIBIASEN,
  TXQPISTRONGPDOWN,
  TXQPIWEAKPUP,
  TXRATE,
  TXSEQUENCE,
  TXSTARTSEQ,
  TXSWING,
  TXSYSCLKSEL,
  TXUSERRDY,
  TXUSRCLK,
  TXUSRCLK2
);

  parameter LOC = "UNPLACED";
  parameter ALIGN_COMMA_DOUBLE = "FALSE";
  parameter [9:0] ALIGN_COMMA_ENABLE = 10'b0001111111;
  parameter integer ALIGN_COMMA_WORD = 1;
  parameter ALIGN_MCOMMA_DET = "TRUE";
  parameter [9:0] ALIGN_MCOMMA_VALUE = 10'b1010000011;
  parameter ALIGN_PCOMMA_DET = "TRUE";
  parameter [9:0] ALIGN_PCOMMA_VALUE = 10'b0101111100;
  parameter CBCC_DATA_SOURCE_SEL = "DECODED";
  parameter CHAN_BOND_KEEP_ALIGN = "FALSE";
  parameter integer CHAN_BOND_MAX_SKEW = 7;
  parameter [9:0] CHAN_BOND_SEQ_1_1 = 10'b0101111100;
  parameter [9:0] CHAN_BOND_SEQ_1_2 = 10'b0000000000;
  parameter [9:0] CHAN_BOND_SEQ_1_3 = 10'b0000000000;
  parameter [9:0] CHAN_BOND_SEQ_1_4 = 10'b0000000000;
  parameter [3:0] CHAN_BOND_SEQ_1_ENABLE = 4'b1111;
  parameter [9:0] CHAN_BOND_SEQ_2_1 = 10'b0100000000;
  parameter [9:0] CHAN_BOND_SEQ_2_2 = 10'b0100000000;
  parameter [9:0] CHAN_BOND_SEQ_2_3 = 10'b0100000000;
  parameter [9:0] CHAN_BOND_SEQ_2_4 = 10'b0100000000;
  parameter [3:0] CHAN_BOND_SEQ_2_ENABLE = 4'b1111;
  parameter CHAN_BOND_SEQ_2_USE = "FALSE";
  parameter integer CHAN_BOND_SEQ_LEN = 1;
  parameter CLK_CORRECT_USE = "TRUE";
  parameter CLK_COR_KEEP_IDLE = "FALSE";
  parameter integer CLK_COR_MAX_LAT = 20;
  parameter integer CLK_COR_MIN_LAT = 18;
  parameter CLK_COR_PRECEDENCE = "TRUE";
  parameter integer CLK_COR_REPEAT_WAIT = 0;
  parameter [9:0] CLK_COR_SEQ_1_1 = 10'b0100011100;
  parameter [9:0] CLK_COR_SEQ_1_2 = 10'b0000000000;
  parameter [9:0] CLK_COR_SEQ_1_3 = 10'b0000000000;
  parameter [9:0] CLK_COR_SEQ_1_4 = 10'b0000000000;
  parameter [3:0] CLK_COR_SEQ_1_ENABLE = 4'b1111;
  parameter [9:0] CLK_COR_SEQ_2_1 = 10'b0100000000;
  parameter [9:0] CLK_COR_SEQ_2_2 = 10'b0100000000;
  parameter [9:0] CLK_COR_SEQ_2_3 = 10'b0100000000;
  parameter [9:0] CLK_COR_SEQ_2_4 = 10'b0100000000;
  parameter [3:0] CLK_COR_SEQ_2_ENABLE = 4'b1111;
  parameter CLK_COR_SEQ_2_USE = "FALSE";
  parameter integer CLK_COR_SEQ_LEN = 1;
  parameter [23:0] CPLL_CFG = 24'hB007D8;
  parameter integer CPLL_FBDIV = 4;
  parameter integer CPLL_FBDIV_45 = 5;
  parameter [23:0] CPLL_INIT_CFG = 24'h00001E;
  parameter [15:0] CPLL_LOCK_CFG = 16'h01E8;
  parameter integer CPLL_REFCLK_DIV = 1;
  parameter integer CPLL_RXOUT_DIV = 2;
  parameter integer CPLL_TXOUT_DIV = 2;
  parameter DEC_MCOMMA_DETECT = "TRUE";
  parameter DEC_PCOMMA_DETECT = "TRUE";
  parameter DEC_VALID_COMMA_ONLY = "TRUE";
  parameter [23:0] DMONITOR_CFG = 24'h000A00;
  parameter [5:0] ES_CONTROL = 6'b000000;
  parameter ES_ERRDET_EN = "FALSE";
  parameter ES_EYE_SCAN_EN = "FALSE";
  parameter [11:0] ES_HORZ_OFFSET = 12'h010;
  parameter [9:0] ES_PMA_CFG = 10'b0000000000;
  parameter [4:0] ES_PRESCALE = 5'b00000;
  parameter [79:0] ES_QUALIFIER = 80'h00000000000000000000;
  parameter [79:0] ES_QUAL_MASK = 80'h00000000000000000000;
  parameter [79:0] ES_SDATA_MASK = 80'h00000000000000000000;
  parameter [8:0] ES_VERT_OFFSET = 9'b000000000;
  parameter [3:0] FTS_DESKEW_SEQ_ENABLE = 4'b1111;
  parameter [3:0] FTS_LANE_DESKEW_CFG = 4'b1111;
  parameter FTS_LANE_DESKEW_EN = "FALSE";
  parameter [2:0] GEARBOX_MODE = 3'b000;
  parameter [1:0] OUTREFCLK_SEL_INV = 2'b11;
  parameter PCS_PCIE_EN = "FALSE";
  parameter [47:0] PCS_RSVD_ATTR = 48'h000000000000;
  parameter [11:0] PD_TRANS_TIME_FROM_P2 = 12'h03C;
  parameter [7:0] PD_TRANS_TIME_NONE_P2 = 8'h19;
  parameter [7:0] PD_TRANS_TIME_TO_P2 = 8'h64;
  parameter [31:0] PMA_RSV = 32'h00000000;
  parameter [15:0] PMA_RSV2 = 16'h0050;
  parameter [1:0] PMA_RSV3 = 2'b00;
  parameter [4:0] RXBUFRESET_TIME = 5'b00001;
  parameter RXBUF_ADDR_MODE = "FULL";
  parameter [3:0] RXBUF_EIDLE_HI_CNT = 4'b1000;
  parameter [3:0] RXBUF_EIDLE_LO_CNT = 4'b0000;
  parameter RXBUF_EN = "TRUE";
  parameter RXBUF_RESET_ON_CB_CHANGE = "TRUE";
  parameter RXBUF_RESET_ON_COMMAALIGN = "FALSE";
  parameter RXBUF_RESET_ON_EIDLE = "TRUE";
  parameter RXBUF_RESET_ON_RATE_CHANGE = "TRUE";
  parameter integer RXBUF_THRESH_OVFLW = 61;
  parameter RXBUF_THRESH_OVRD = "FALSE";
  parameter integer RXBUF_THRESH_UNDFLW = 4;
  parameter [4:0] RXCDRFREQRESET_TIME = 5'b00001;
  parameter [4:0] RXCDRPHRESET_TIME = 5'b00001;
  parameter [71:0] RXCDR_CFG = 72'h1107FE406001080000;
  parameter [0:0] RXCDR_FR_RESET_ON_EIDLE = 1'b0;
  parameter [0:0] RXCDR_HOLD_DURING_EIDLE = 1'b0;
  parameter [5:0] RXCDR_LOCK_CFG = 6'b001001;
  parameter [0:0] RXCDR_PH_RESET_ON_EIDLE = 1'b0;
  parameter [6:0] RXDFELPMRESET_TIME = 7'b0001111;
  parameter [15:0] RXDLY_CFG = 16'h0010;
  parameter [8:0] RXDLY_LCFG = 9'h020;
  parameter [15:0] RXDLY_TAP_CFG = 16'h0000;
  parameter RXGEARBOX_EN = "FALSE";
  parameter [4:0] RXISCANRESET_TIME = 5'b00001;
  parameter [13:0] RXLPM_HF_CFG = 14'b00001111110000;
  parameter [13:0] RXLPM_LF_CFG = 14'b00001111110000;
  parameter [6:0] RXOOB_CFG = 7'b0000110;
  parameter [4:0] RXPCSRESET_TIME = 5'b00001;
  parameter [23:0] RXPHDLY_CFG = 24'h084000;
  parameter [23:0] RXPH_CFG = 24'h000000;
  parameter [4:0] RXPH_MONITOR_SEL = 5'b00000;
  parameter [4:0] RXPMARESET_TIME = 5'b00011;
  parameter [0:0] RXPRBS_ERR_LOOPBACK = 1'b0;
  parameter integer RXSLIDE_AUTO_WAIT = 5;
  parameter RXSLIDE_MODE = "OFF";
  parameter [11:0] RX_BIAS_CFG = 12'b000000000000;
  parameter [5:0] RX_BUFFER_CFG = 6'b000000;
  parameter integer RX_CLK25_DIV = 7;
  parameter [0:0] RX_CLKMUX_PD = 1'b0;
  parameter [1:0] RX_CM_SEL = 2'b11;
  parameter [2:0] RX_CM_TRIM = 3'b100;
  parameter integer RX_DATA_WIDTH = 20;
  parameter [5:0] RX_DDI_SEL = 6'b000000;
  parameter [11:0] RX_DEBUG_CFG = 12'b000000000000;
  parameter RX_DEFER_RESET_BUF_EN = "TRUE";
  parameter [22:0] RX_DFE_GAIN_CFG = 23'h181C0F;
  parameter [11:0] RX_DFE_H2_CFG = 12'b000111100000;
  parameter [11:0] RX_DFE_H3_CFG = 12'b000111100000;
  parameter [10:0] RX_DFE_H4_CFG = 11'b00011110000;
  parameter [10:0] RX_DFE_H5_CFG = 11'b00011110000;
  parameter [12:0] RX_DFE_KL_CFG = 13'b0001111110000;
  parameter [15:0] RX_DFE_LPM_CFG = 16'h0000;
  parameter [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE = 1'b0;
  parameter [16:0] RX_DFE_UT_CFG = 17'b00011111100000000;
  parameter [16:0] RX_DFE_VP_CFG = 17'b00011111100000000;
  parameter [12:0] RX_DFE_XYD_CFG = 13'b0001100010000;
  parameter RX_DISPERR_SEQ_MATCH = "TRUE";
  parameter integer RX_INT_DATAWIDTH = 0;
  parameter [12:0] RX_OS_CFG = 13'b0001111110000;
  parameter integer RX_SIG_VALID_DLY = 10;
  parameter RX_XCLK_SEL = "RXREC";
  parameter integer SAS_MAX_COM = 64;
  parameter integer SAS_MIN_COM = 36;
  parameter [3:0] SATA_BURST_SEQ_LEN = 4'b1111;
  parameter [2:0] SATA_BURST_VAL = 3'b100;
  parameter SATA_CPLL_CFG = "VCO_3000MHZ";
  parameter [2:0] SATA_EIDLE_VAL = 3'b100;
  parameter integer SATA_MAX_BURST = 8;
  parameter integer SATA_MAX_INIT = 21;
  parameter integer SATA_MAX_WAKE = 7;
  parameter integer SATA_MIN_BURST = 4;
  parameter integer SATA_MIN_INIT = 12;
  parameter integer SATA_MIN_WAKE = 4;
  parameter SHOW_REALIGN_COMMA = "TRUE";
  parameter [2:0] SIM_CPLLREFCLK_SEL = 3'b001;
  parameter SIM_RECEIVER_DETECT_PASS = "TRUE";
  parameter SIM_RESET_SPEEDUP = "TRUE";
  parameter SIM_TX_EIDLE_DRIVE_LEVEL = "X";
  parameter SIM_VERSION = "1.0";
  parameter [4:0] TERM_RCAL_CFG = 5'b10000;
  parameter [0:0] TERM_RCAL_OVRD = 1'b0;
  parameter [7:0] TRANS_TIME_RATE = 8'h0E;
  parameter [31:0] TST_RSV = 32'h00000000;
  parameter TXBUF_EN = "TRUE";
  parameter TXBUF_RESET_ON_RATE_CHANGE = "FALSE";
  parameter [15:0] TXDLY_CFG = 16'h0010;
  parameter [8:0] TXDLY_LCFG = 9'h020;
  parameter [15:0] TXDLY_TAP_CFG = 16'h0000;
  parameter TXGEARBOX_EN = "FALSE";
  parameter [4:0] TXPCSRESET_TIME = 5'b00001;
  parameter [23:0] TXPHDLY_CFG = 24'h084000;
  parameter [15:0] TXPH_CFG = 16'h0400;
  parameter [4:0] TXPH_MONITOR_SEL = 5'b00000;
  parameter [4:0] TXPMARESET_TIME = 5'b00001;
  parameter integer TX_CLK25_DIV = 7;
  parameter [0:0] TX_CLKMUX_PD = 1'b0;
  parameter integer TX_DATA_WIDTH = 20;
  parameter [4:0] TX_DEEMPH0 = 5'b00000;
  parameter [4:0] TX_DEEMPH1 = 5'b00000;
  parameter TX_DRIVE_MODE = "DIRECT";
  parameter [2:0] TX_EIDLE_ASSERT_DELAY = 3'b110;
  parameter [2:0] TX_EIDLE_DEASSERT_DELAY = 3'b100;
  parameter integer TX_INT_DATAWIDTH = 0;
  parameter TX_LOOPBACK_DRIVE_HIZ = "FALSE";
  parameter [0:0] TX_MAINCURSOR_SEL = 1'b0;
  parameter [6:0] TX_MARGIN_FULL_0 = 7'b1001110;
  parameter [6:0] TX_MARGIN_FULL_1 = 7'b1001001;
  parameter [6:0] TX_MARGIN_FULL_2 = 7'b1000101;
  parameter [6:0] TX_MARGIN_FULL_3 = 7'b1000010;
  parameter [6:0] TX_MARGIN_FULL_4 = 7'b1000000;
  parameter [6:0] TX_MARGIN_LOW_0 = 7'b1000110;
  parameter [6:0] TX_MARGIN_LOW_1 = 7'b1000100;
  parameter [6:0] TX_MARGIN_LOW_2 = 7'b1000010;
  parameter [6:0] TX_MARGIN_LOW_3 = 7'b1000000;
  parameter [6:0] TX_MARGIN_LOW_4 = 7'b1000000;
  parameter [0:0] TX_PREDRIVER_MODE = 1'b0;
  parameter [0:0] TX_QPI_STATUS_EN = 1'b0;
  parameter [13:0] TX_RXDETECT_CFG = 14'h1832;
  parameter [2:0] TX_RXDETECT_REF = 3'b100;
  parameter TX_XCLK_SEL = "TXUSR";
  parameter [0:0] UCODEER_CLR = 1'b0;
  
  localparam in_delay = 0;
  localparam out_delay = 0;
  localparam INCLK_DELAY = 0;
  localparam OUTCLK_DELAY = 0;

  output CPLLFBCLKLOST;
  output CPLLLOCK;
  output CPLLREFCLKLOST;
  output DRPRDY;
  output EYESCANDATAERROR;
  output GTREFCLKMONITOR;
  output GTXTXN;
  output GTXTXP;
  output PHYSTATUS;
  output RXBYTEISALIGNED;
  output RXBYTEREALIGN;
  output RXCDRLOCK;
  output RXCHANBONDSEQ;
  output RXCHANISALIGNED;
  output RXCHANREALIGN;
  output RXCOMINITDET;
  output RXCOMMADET;
  output RXCOMSASDET;
  output RXCOMWAKEDET;
  output RXDATAVALID;
  output RXDLYSRESETDONE;
  output RXELECIDLE;
  output RXHEADERVALID;
  output RXOUTCLK;
  output RXOUTCLKFABRIC;
  output RXOUTCLKPCS;
  output RXPHALIGNDONE;
  output RXPRBSERR;
  output RXQPISENN;
  output RXQPISENP;
  output RXRATEDONE;
  output RXRESETDONE;
  output RXSTARTOFSEQ;
  output RXVALID;
  output TXCOMFINISH;
  output TXDLYSRESETDONE;
  output TXGEARBOXREADY;
  output TXOUTCLK;
  output TXOUTCLKFABRIC;
  output TXOUTCLKPCS;
  output TXPHALIGNDONE;
  output TXPHINITDONE;
  output TXQPISENN;
  output TXQPISENP;
  output TXRATEDONE;
  output TXRESETDONE;
  output [15:0] DRPDO;
  output [15:0] PCSRSVDOUT;
  output [1:0] RXCLKCORCNT;
  output [1:0] TXBUFSTATUS;
  output [2:0] RXBUFSTATUS;
  output [2:0] RXHEADER;
  output [2:0] RXSTATUS;
  output [4:0] RXCHBONDO;
  output [4:0] RXPHMONITOR;
  output [4:0] RXPHSLIPMONITOR;
  output [63:0] RXDATA;
  output [6:0] RXMONITOROUT;
  output [7:0] DMONITOROUT;
  output [7:0] RXCHARISCOMMA;
  output [7:0] RXCHARISK;
  output [7:0] RXDISPERR;
  output [7:0] RXNOTINTABLE;
  output [9:0] TSTOUT;

  input CFGRESET;
  input CPLLLOCKDETCLK;
  input CPLLLOCKEN;
  input CPLLPD;
  input CPLLRESET;
  input DRPCLK;
  input DRPEN;
  input DRPWE;
  input EYESCANMODE;
  input EYESCANRESET;
  input EYESCANTRIGGER;
  input GTGREFCLK;
  input GTNORTHREFCLK0;
  input GTNORTHREFCLK1;
  input GTREFCLK0;
  input GTREFCLK1;
  input GTRESETSEL;
  input GTRXRESET;
  input GTSOUTHREFCLK0;
  input GTSOUTHREFCLK1;
  input GTTXRESET;
  input GTXRXN;
  input GTXRXP;
  input QPLLCLK;
  input QPLLREFCLK;
  input RESETOVRD;
  input RX8B10BEN;
  input RXBUFRESET;
  input RXCDRFREQRESET;
  input RXCDRHOLD;
  input RXCDROVRDEN;
  input RXCDRRESET;
  input RXCDRRESETRSV;
  input RXCHBONDEN;
  input RXCHBONDMASTER;
  input RXCHBONDSLAVE;
  input RXCOMMADETEN;
  input RXDDIEN;
  input RXDFEAGCHOLD;
  input RXDFEAGCOVRDEN;
  input RXDFECM1EN;
  input RXDFELFHOLD;
  input RXDFELFOVRDEN;
  input RXDFELPMRESET;
  input RXDFETAP2HOLD;
  input RXDFETAP2OVRDEN;
  input RXDFETAP3HOLD;
  input RXDFETAP3OVRDEN;
  input RXDFETAP4HOLD;
  input RXDFETAP4OVRDEN;
  input RXDFETAP5HOLD;
  input RXDFETAP5OVRDEN;
  input RXDFEUTHOLD;
  input RXDFEUTOVRDEN;
  input RXDFEVPHOLD;
  input RXDFEVPOVRDEN;
  input RXDFEVSEN;
  input RXDFEXYDEN;
  input RXDFEXYDHOLD;
  input RXDFEXYDOVRDEN;
  input RXDLYBYPASS;
  input RXDLYEN;
  input RXDLYOVRDEN;
  input RXDLYSRESET;
  input RXGEARBOXSLIP;
  input RXLPMEN;
  input RXLPMHFHOLD;
  input RXLPMHFOVRDEN;
  input RXLPMLFHOLD;
  input RXLPMLFKLOVRDEN;
  input RXMCOMMAALIGNEN;
  input RXOOBRESET;
  input RXOSHOLD;
  input RXOSOVRDEN;
  input RXPCOMMAALIGNEN;
  input RXPCSRESET;
  input RXPHALIGN;
  input RXPHALIGNEN;
  input RXPHDLYPD;
  input RXPHDLYRESET;
  input RXPHOVRDEN;
  input RXPMARESET;
  input RXPOLARITY;
  input RXPRBSCNTRESET;
  input RXQPIEN;
  input RXSLIDE;
  input RXUSERRDY;
  input RXUSRCLK2;
  input RXUSRCLK;
  input SETERRSTATUS;
  input TX8B10BEN;
  input TXCOMINIT;
  input TXCOMSAS;
  input TXCOMWAKE;
  input TXDEEMPH;
  input TXDETECTRX;
  input TXDIFFPD;
  input TXDLYBYPASS;
  input TXDLYEN;
  input TXDLYHOLD;
  input TXDLYOVRDEN;
  input TXDLYSRESET;
  input TXDLYUPDOWN;
  input TXELECIDLE;
  input TXINHIBIT;
  input TXPCSRESET;
  input TXPDELECIDLEMODE;
  input TXPHALIGN;
  input TXPHALIGNEN;
  input TXPHDLYPD;
  input TXPHDLYRESET;
  input TXPHDLYTSTCLK;
  input TXPHINIT;
  input TXPHOVRDEN;
  input TXPISOPD;
  input TXPMARESET;
  input TXPOLARITY;
  input TXPOSTCURSORINV;
  input TXPRBSFORCEERR;
  input TXPRECURSORINV;
  input TXQPIBIASEN;
  input TXQPISTRONGPDOWN;
  input TXQPIWEAKPUP;
  input TXSTARTSEQ;
  input TXSWING;
  input TXUSERRDY;
  input TXUSRCLK2;
  input TXUSRCLK;
  input [15:0] DRPDI;
  input [15:0] GTRSVD;
  input [15:0] PCSRSVDIN;
  input [19:0] TSTIN;
  input [1:0] RXELECIDLEMODE;
  input [1:0] RXMONITORSEL;
  input [1:0] RXPD;
  input [1:0] RXSYSCLKSEL;
  input [1:0] TXPD;
  input [1:0] TXSYSCLKSEL;
  input [2:0] CPLLREFCLKSEL;
  input [2:0] LOOPBACK;
  input [2:0] RXCHBONDLEVEL;
  input [2:0] RXOUTCLKSEL;
  input [2:0] RXPRBSSEL;
  input [2:0] RXRATE;
  input [2:0] TXBUFDIFFCTRL;
  input [2:0] TXHEADER;
  input [2:0] TXMARGIN;
  input [2:0] TXOUTCLKSEL;
  input [2:0] TXPRBSSEL;
  input [2:0] TXRATE;
  input [3:0] CLKRSVD;
  input [3:0] TXDIFFCTRL;
  input [4:0] PCSRSVDIN2;
  input [4:0] PMARSVDIN2;
  input [4:0] PMARSVDIN;
  input [4:0] RXCHBONDI;
  input [4:0] TXPOSTCURSOR;
  input [4:0] TXPRECURSOR;
  input [63:0] TXDATA;
  input [6:0] TXMAINCURSOR;
  input [6:0] TXSEQUENCE;
  input [7:0] TX8B10BBYPASS;
  input [7:0] TXCHARDISPMODE;
  input [7:0] TXCHARDISPVAL;
  input [7:0] TXCHARISK;
  input [8:0] DRPADDR;

  reg SIM_RECEIVER_DETECT_PASS_BINARY;
  reg SIM_RESET_SPEEDUP_BINARY;
  reg SIM_TX_EIDLE_DRIVE_LEVEL_BINARY;
  reg SIM_VERSION_BINARY;
  reg [0:0] ALIGN_COMMA_DOUBLE_BINARY;
  reg [0:0] ALIGN_MCOMMA_DET_BINARY;
  reg [0:0] ALIGN_PCOMMA_DET_BINARY;
  reg [0:0] CBCC_DATA_SOURCE_SEL_BINARY;
  reg [0:0] CHAN_BOND_KEEP_ALIGN_BINARY;
  reg [0:0] CHAN_BOND_SEQ_2_USE_BINARY;
  reg [0:0] CLK_CORRECT_USE_BINARY;
  reg [0:0] CLK_COR_KEEP_IDLE_BINARY;
  reg [0:0] CLK_COR_PRECEDENCE_BINARY;
  reg [0:0] CLK_COR_SEQ_2_USE_BINARY;
  reg [0:0] CPLL_FBDIV_45_BINARY;
  reg [0:0] DEC_MCOMMA_DETECT_BINARY;
  reg [0:0] DEC_PCOMMA_DETECT_BINARY;
  reg [0:0] DEC_VALID_COMMA_ONLY_BINARY;
  reg [0:0] ES_ERRDET_EN_BINARY;
  reg [0:0] ES_EYE_SCAN_EN_BINARY;
  reg [0:0] FTS_LANE_DESKEW_EN_BINARY;
  reg [0:0] PCS_PCIE_EN_BINARY;
  reg [0:0] RXBUF_ADDR_MODE_BINARY;
  reg [0:0] RXBUF_EN_BINARY;
  reg [0:0] RXBUF_RESET_ON_CB_CHANGE_BINARY;
  reg [0:0] RXBUF_RESET_ON_COMMAALIGN_BINARY;
  reg [0:0] RXBUF_RESET_ON_EIDLE_BINARY;
  reg [0:0] RXBUF_RESET_ON_RATE_CHANGE_BINARY;
  reg [0:0] RXBUF_THRESH_OVRD_BINARY;
  reg [0:0] RXCDR_FR_RESET_ON_EIDLE_BINARY;
  reg [0:0] RXCDR_HOLD_DURING_EIDLE_BINARY;
  reg [0:0] RXCDR_PH_RESET_ON_EIDLE_BINARY;
  reg [0:0] RXGEARBOX_EN_BINARY;
  reg [0:0] RXPRBS_ERR_LOOPBACK_BINARY;
  reg [0:0] RX_CLKMUX_PD_BINARY;
  reg [0:0] RX_DEFER_RESET_BUF_EN_BINARY;
  reg [0:0] RX_DFE_LPM_HOLD_DURING_EIDLE_BINARY;
  reg [0:0] RX_DISPERR_SEQ_MATCH_BINARY;
  reg [0:0] RX_INT_DATAWIDTH_BINARY;
  reg [0:0] RX_XCLK_SEL_BINARY;
  reg [0:0] SHOW_REALIGN_COMMA_BINARY;
  reg [0:0] TERM_RCAL_OVRD_BINARY;
  reg [0:0] TXBUF_EN_BINARY;
  reg [0:0] TXBUF_RESET_ON_RATE_CHANGE_BINARY;
  reg [0:0] TXGEARBOX_EN_BINARY;
  reg [0:0] TX_CLKMUX_PD_BINARY;
  reg [0:0] TX_INT_DATAWIDTH_BINARY;
  reg [0:0] TX_LOOPBACK_DRIVE_HIZ_BINARY;
  reg [0:0] TX_MAINCURSOR_SEL_BINARY;
  reg [0:0] TX_PREDRIVER_MODE_BINARY;
  reg [0:0] TX_QPI_STATUS_EN_BINARY;
  reg [0:0] TX_XCLK_SEL_BINARY;
  reg [0:0] UCODEER_CLR_BINARY;
  reg [10:0] RX_DFE_H4_CFG_BINARY;
  reg [10:0] RX_DFE_H5_CFG_BINARY;
  reg [11:0] RX_BIAS_CFG_BINARY;
  reg [11:0] RX_DEBUG_CFG_BINARY;
  reg [11:0] RX_DFE_H2_CFG_BINARY;
  reg [11:0] RX_DFE_H3_CFG_BINARY;
  reg [12:0] RX_DFE_KL_CFG_BINARY;
  reg [12:0] RX_DFE_XYD_CFG_BINARY;
  reg [12:0] RX_OS_CFG_BINARY;
  reg [13:0] RXLPM_HF_CFG_BINARY;
  reg [13:0] RXLPM_LF_CFG_BINARY;
  reg [16:0] RX_DFE_UT_CFG_BINARY;
  reg [16:0] RX_DFE_VP_CFG_BINARY;
  reg [1:0] CHAN_BOND_SEQ_LEN_BINARY;
  reg [1:0] CLK_COR_SEQ_LEN_BINARY;
  reg [1:0] OUTREFCLK_SEL_INV_BINARY;
  reg [1:0] PMA_RSV3_BINARY;
  reg [1:0] RXSLIDE_MODE_BINARY;
  reg [1:0] RX_CM_SEL_BINARY;
  reg [1:0] SATA_CPLL_CFG_BINARY;
  reg [2:0] ALIGN_COMMA_WORD_BINARY;
  reg [2:0] CPLL_RXOUT_DIV_BINARY;
  reg [2:0] CPLL_TXOUT_DIV_BINARY;
  reg [2:0] GEARBOX_MODE_BINARY;
  reg [2:0] RX_CM_TRIM_BINARY;
  reg [2:0] RX_DATA_WIDTH_BINARY;
  reg [2:0] SATA_BURST_VAL_BINARY;
  reg [2:0] SATA_EIDLE_VAL_BINARY;
  reg [2:0] SIM_CPLLREFCLK_SEL_BINARY;
  reg [2:0] TX_DATA_WIDTH_BINARY;
  reg [2:0] TX_EIDLE_ASSERT_DELAY_BINARY;
  reg [2:0] TX_EIDLE_DEASSERT_DELAY_BINARY;
  reg [2:0] TX_RXDETECT_REF_BINARY;
  reg [3:0] CHAN_BOND_MAX_SKEW_BINARY;
  reg [3:0] CHAN_BOND_SEQ_1_ENABLE_BINARY;
  reg [3:0] CHAN_BOND_SEQ_2_ENABLE_BINARY;
  reg [3:0] CLK_COR_SEQ_1_ENABLE_BINARY;
  reg [3:0] CLK_COR_SEQ_2_ENABLE_BINARY;
  reg [3:0] FTS_DESKEW_SEQ_ENABLE_BINARY;
  reg [3:0] FTS_LANE_DESKEW_CFG_BINARY;
  reg [3:0] RXBUF_EIDLE_HI_CNT_BINARY;
  reg [3:0] RXBUF_EIDLE_LO_CNT_BINARY;
  reg [3:0] RXSLIDE_AUTO_WAIT_BINARY;
  reg [3:0] SATA_BURST_SEQ_LEN_BINARY;
  reg [4:0] CLK_COR_REPEAT_WAIT_BINARY;
  reg [4:0] CPLL_REFCLK_DIV_BINARY;
  reg [4:0] ES_PRESCALE_BINARY;
  reg [4:0] RXBUFRESET_TIME_BINARY;
  reg [4:0] RXCDRFREQRESET_TIME_BINARY;
  reg [4:0] RXCDRPHRESET_TIME_BINARY;
  reg [4:0] RXISCANRESET_TIME_BINARY;
  reg [4:0] RXPCSRESET_TIME_BINARY;
  reg [4:0] RXPH_MONITOR_SEL_BINARY;
  reg [4:0] RXPMARESET_TIME_BINARY;
  reg [4:0] RX_CLK25_DIV_BINARY;
  reg [4:0] RX_SIG_VALID_DLY_BINARY;
  reg [4:0] TERM_RCAL_CFG_BINARY;
  reg [4:0] TXPCSRESET_TIME_BINARY;
  reg [4:0] TXPH_MONITOR_SEL_BINARY;
  reg [4:0] TXPMARESET_TIME_BINARY;
  reg [4:0] TX_CLK25_DIV_BINARY;
  reg [4:0] TX_DEEMPH0_BINARY;
  reg [4:0] TX_DEEMPH1_BINARY;
  reg [4:0] TX_DRIVE_MODE_BINARY;
  reg [5:0] CLK_COR_MAX_LAT_BINARY;
  reg [5:0] CLK_COR_MIN_LAT_BINARY;
  reg [5:0] ES_CONTROL_BINARY;
  reg [5:0] RXBUF_THRESH_OVFLW_BINARY;
  reg [5:0] RXBUF_THRESH_UNDFLW_BINARY;
  reg [5:0] RXCDR_LOCK_CFG_BINARY;
  reg [5:0] RX_BUFFER_CFG_BINARY;
  reg [5:0] RX_DDI_SEL_BINARY;
  reg [5:0] SAS_MIN_COM_BINARY;
  reg [5:0] SATA_MAX_BURST_BINARY;
  reg [5:0] SATA_MAX_INIT_BINARY;
  reg [5:0] SATA_MAX_WAKE_BINARY;
  reg [5:0] SATA_MIN_BURST_BINARY;
  reg [5:0] SATA_MIN_INIT_BINARY;
  reg [5:0] SATA_MIN_WAKE_BINARY;
  reg [6:0] CPLL_FBDIV_BINARY;
  reg [6:0] RXDFELPMRESET_TIME_BINARY;
  reg [6:0] RXOOB_CFG_BINARY;
  reg [6:0] SAS_MAX_COM_BINARY;
  reg [6:0] TX_MARGIN_FULL_0_BINARY;
  reg [6:0] TX_MARGIN_FULL_1_BINARY;
  reg [6:0] TX_MARGIN_FULL_2_BINARY;
  reg [6:0] TX_MARGIN_FULL_3_BINARY;
  reg [6:0] TX_MARGIN_FULL_4_BINARY;
  reg [6:0] TX_MARGIN_LOW_0_BINARY;
  reg [6:0] TX_MARGIN_LOW_1_BINARY;
  reg [6:0] TX_MARGIN_LOW_2_BINARY;
  reg [6:0] TX_MARGIN_LOW_3_BINARY;
  reg [6:0] TX_MARGIN_LOW_4_BINARY;
  reg [8:0] ES_VERT_OFFSET_BINARY;
  reg [9:0] ALIGN_COMMA_ENABLE_BINARY;
  reg [9:0] ALIGN_MCOMMA_VALUE_BINARY;
  reg [9:0] ALIGN_PCOMMA_VALUE_BINARY;
  reg [9:0] CHAN_BOND_SEQ_1_1_BINARY;
  reg [9:0] CHAN_BOND_SEQ_1_2_BINARY;
  reg [9:0] CHAN_BOND_SEQ_1_3_BINARY;
  reg [9:0] CHAN_BOND_SEQ_1_4_BINARY;
  reg [9:0] CHAN_BOND_SEQ_2_1_BINARY;
  reg [9:0] CHAN_BOND_SEQ_2_2_BINARY;
  reg [9:0] CHAN_BOND_SEQ_2_3_BINARY;
  reg [9:0] CHAN_BOND_SEQ_2_4_BINARY;
  reg [9:0] CLK_COR_SEQ_1_1_BINARY;
  reg [9:0] CLK_COR_SEQ_1_2_BINARY;
  reg [9:0] CLK_COR_SEQ_1_3_BINARY;
  reg [9:0] CLK_COR_SEQ_1_4_BINARY;
  reg [9:0] CLK_COR_SEQ_2_1_BINARY;
  reg [9:0] CLK_COR_SEQ_2_2_BINARY;
  reg [9:0] CLK_COR_SEQ_2_3_BINARY;
  reg [9:0] CLK_COR_SEQ_2_4_BINARY;
  reg [9:0] ES_PMA_CFG_BINARY;

  tri0 GSR = glbl.GSR;
  reg notifier;

  wire CPLLFBCLKLOST_OUT;
  wire CPLLLOCK_OUT;
  wire CPLLREFCLKLOST_OUT;
  wire DRPRDY_OUT;
  wire EYESCANDATAERROR_OUT;
  wire GTREFCLKMONITOR_OUT;
  wire GTXTXN_OUT;
  wire GTXTXP_OUT;
  wire PHYSTATUS_OUT;
  wire RXBYTEISALIGNED_OUT;
  wire RXBYTEREALIGN_OUT;
  wire RXCDRLOCK_OUT;
  wire RXCHANBONDSEQ_OUT;
  wire RXCHANISALIGNED_OUT;
  wire RXCHANREALIGN_OUT;
  wire RXCOMINITDET_OUT;
  wire RXCOMMADET_OUT;
  wire RXCOMSASDET_OUT;
  wire RXCOMWAKEDET_OUT;
  wire RXDATAVALID_OUT;
  wire RXDLYSRESETDONE_OUT;
  wire RXELECIDLE_OUT;
  wire RXHEADERVALID_OUT;
  wire RXOUTCLKFABRIC_OUT;
  wire RXOUTCLKPCS_OUT;
  wire RXOUTCLK_OUT;
  wire RXPHALIGNDONE_OUT;
  wire RXPRBSERR_OUT;
  wire RXQPISENN_OUT;
  wire RXQPISENP_OUT;
  wire RXRATEDONE_OUT;
  wire RXRESETDONE_OUT;
  wire RXSTARTOFSEQ_OUT;
  wire RXVALID_OUT;
  wire TXCOMFINISH_OUT;
  wire TXDLYSRESETDONE_OUT;
  wire TXGEARBOXREADY_OUT;
  wire TXOUTCLKFABRIC_OUT;
  wire TXOUTCLKPCS_OUT;
  wire TXOUTCLK_OUT;
  wire TXPHALIGNDONE_OUT;
  wire TXPHINITDONE_OUT;
  wire TXQPISENN_OUT;
  wire TXQPISENP_OUT;
  wire TXRATEDONE_OUT;
  wire TXRESETDONE_OUT;
  wire [15:0] DRPDO_OUT;
  wire [15:0] PCSRSVDOUT_OUT;
  wire [1:0] RXCLKCORCNT_OUT;
  wire [1:0] TXBUFSTATUS_OUT;
  wire [2:0] RXBUFSTATUS_OUT;
  wire [2:0] RXHEADER_OUT;
  wire [2:0] RXSTATUS_OUT;
  wire [4:0] RXCHBONDO_OUT;
  wire [4:0] RXPHMONITOR_OUT;
  wire [4:0] RXPHSLIPMONITOR_OUT;
  wire [63:0] RXDATA_OUT;
  wire [6:0] RXMONITOROUT_OUT;
  wire [7:0] DMONITOROUT_OUT;
  wire [7:0] RXCHARISCOMMA_OUT;
  wire [7:0] RXCHARISK_OUT;
  wire [7:0] RXDISPERR_OUT;
  wire [7:0] RXNOTINTABLE_OUT;
  wire [9:0] TSTOUT_OUT;

  wire CFGRESET_IN;
  wire CPLLLOCKDETCLK_IN;
  wire CPLLLOCKEN_IN;
  wire CPLLPD_IN;
  wire CPLLRESET_IN;
  wire DRPCLK_IN;
  wire DRPEN_IN;
  wire DRPWE_IN;
  wire EYESCANMODE_IN;
  wire EYESCANRESET_IN;
  wire EYESCANTRIGGER_IN;
  wire GTGREFCLK_IN;
  wire GTNORTHREFCLK0_IN;
  wire GTNORTHREFCLK1_IN;
  wire GTREFCLK0_IN;
  wire GTREFCLK1_IN;
  wire GTRESETSEL_IN;
  wire GTRXRESET_IN;
  wire GTSOUTHREFCLK0_IN;
  wire GTSOUTHREFCLK1_IN;
  wire GTTXRESET_IN;
  wire GTXRXN_IN;
  wire GTXRXP_IN;
  wire QPLLCLK_IN;
  wire QPLLREFCLK_IN;
  wire RESETOVRD_IN;
  wire RX8B10BEN_IN;
  wire RXBUFRESET_IN;
  wire RXCDRFREQRESET_IN;
  wire RXCDRHOLD_IN;
  wire RXCDROVRDEN_IN;
  wire RXCDRRESETRSV_IN;
  wire RXCDRRESET_IN;
  wire RXCHBONDEN_IN;
  wire RXCHBONDMASTER_IN;
  wire RXCHBONDSLAVE_IN;
  wire RXCOMMADETEN_IN;
  wire RXDDIEN_IN;
  wire RXDFEAGCHOLD_IN;
  wire RXDFEAGCOVRDEN_IN;
  wire RXDFECM1EN_IN;
  wire RXDFELFHOLD_IN;
  wire RXDFELFOVRDEN_IN;
  wire RXDFELPMRESET_IN;
  wire RXDFETAP2HOLD_IN;
  wire RXDFETAP2OVRDEN_IN;
  wire RXDFETAP3HOLD_IN;
  wire RXDFETAP3OVRDEN_IN;
  wire RXDFETAP4HOLD_IN;
  wire RXDFETAP4OVRDEN_IN;
  wire RXDFETAP5HOLD_IN;
  wire RXDFETAP5OVRDEN_IN;
  wire RXDFEUTHOLD_IN;
  wire RXDFEUTOVRDEN_IN;
  wire RXDFEVPHOLD_IN;
  wire RXDFEVPOVRDEN_IN;
  wire RXDFEVSEN_IN;
  wire RXDFEXYDEN_IN;
  wire RXDFEXYDHOLD_IN;
  wire RXDFEXYDOVRDEN_IN;
  wire RXDLYBYPASS_IN;
  wire RXDLYEN_IN;
  wire RXDLYOVRDEN_IN;
  wire RXDLYSRESET_IN;
  wire RXGEARBOXSLIP_IN;
  wire RXLPMEN_IN;
  wire RXLPMHFHOLD_IN;
  wire RXLPMHFOVRDEN_IN;
  wire RXLPMLFHOLD_IN;
  wire RXLPMLFKLOVRDEN_IN;
  wire RXMCOMMAALIGNEN_IN;
  wire RXOOBRESET_IN;
  wire RXOSHOLD_IN;
  wire RXOSOVRDEN_IN;
  wire RXPCOMMAALIGNEN_IN;
  wire RXPCSRESET_IN;
  wire RXPHALIGNEN_IN;
  wire RXPHALIGN_IN;
  wire RXPHDLYPD_IN;
  wire RXPHDLYRESET_IN;
  wire RXPHOVRDEN_IN;
  wire RXPMARESET_IN;
  wire RXPOLARITY_IN;
  wire RXPRBSCNTRESET_IN;
  wire RXQPIEN_IN;
  wire RXSLIDE_IN;
  wire RXUSERRDY_IN;
  wire RXUSRCLK2_IN;
  wire RXUSRCLK_IN;
  wire SETERRSTATUS_IN;
  wire TX8B10BEN_IN;
  wire TXCOMINIT_IN;
  wire TXCOMSAS_IN;
  wire TXCOMWAKE_IN;
  wire TXDEEMPH_IN;
  wire TXDETECTRX_IN;
  wire TXDIFFPD_IN;
  wire TXDLYBYPASS_IN;
  wire TXDLYEN_IN;
  wire TXDLYHOLD_IN;
  wire TXDLYOVRDEN_IN;
  wire TXDLYSRESET_IN;
  wire TXDLYUPDOWN_IN;
  wire TXELECIDLE_IN;
  wire TXINHIBIT_IN;
  wire TXPCSRESET_IN;
  wire TXPDELECIDLEMODE_IN;
  wire TXPHALIGNEN_IN;
  wire TXPHALIGN_IN;
  wire TXPHDLYPD_IN;
  wire TXPHDLYRESET_IN;
  wire TXPHDLYTSTCLK_IN;
  wire TXPHINIT_IN;
  wire TXPHOVRDEN_IN;
  wire TXPISOPD_IN;
  wire TXPMARESET_IN;
  wire TXPOLARITY_IN;
  wire TXPOSTCURSORINV_IN;
  wire TXPRBSFORCEERR_IN;
  wire TXPRECURSORINV_IN;
  wire TXQPIBIASEN_IN;
  wire TXQPISTRONGPDOWN_IN;
  wire TXQPIWEAKPUP_IN;
  wire TXSTARTSEQ_IN;
  wire TXSWING_IN;
  wire TXUSERRDY_IN;
  wire TXUSRCLK2_IN;
  wire TXUSRCLK_IN;
  wire [15:0] DRPDI_IN;
  wire [15:0] GTRSVD_IN;
  wire [15:0] PCSRSVDIN_IN;
  wire [19:0] TSTIN_IN;
  wire [1:0] RXELECIDLEMODE_IN;
  wire [1:0] RXMONITORSEL_IN;
  wire [1:0] RXPD_IN;
  wire [1:0] RXSYSCLKSEL_IN;
  wire [1:0] TXPD_IN;
  wire [1:0] TXSYSCLKSEL_IN;
  wire [2:0] CPLLREFCLKSEL_IN;
  wire [2:0] LOOPBACK_IN;
  wire [2:0] RXCHBONDLEVEL_IN;
  wire [2:0] RXOUTCLKSEL_IN;
  wire [2:0] RXPRBSSEL_IN;
  wire [2:0] RXRATE_IN;
  wire [2:0] TXBUFDIFFCTRL_IN;
  wire [2:0] TXHEADER_IN;
  wire [2:0] TXMARGIN_IN;
  wire [2:0] TXOUTCLKSEL_IN;
  wire [2:0] TXPRBSSEL_IN;
  wire [2:0] TXRATE_IN;
  wire [3:0] CLKRSVD_IN;
  wire [3:0] TXDIFFCTRL_IN;
  wire [4:0] PCSRSVDIN2_IN;
  wire [4:0] PMARSVDIN2_IN;
  wire [4:0] PMARSVDIN_IN;
  wire [4:0] RXCHBONDI_IN;
  wire [4:0] TXPOSTCURSOR_IN;
  wire [4:0] TXPRECURSOR_IN;
  wire [63:0] TXDATA_IN;
  wire [6:0] TXMAINCURSOR_IN;
  wire [6:0] TXSEQUENCE_IN;
  wire [7:0] TX8B10BBYPASS_IN;
  wire [7:0] TXCHARDISPMODE_IN;
  wire [7:0] TXCHARDISPVAL_IN;
  wire [7:0] TXCHARISK_IN;
  wire [8:0] DRPADDR_IN;

  wire CFGRESET_INDELAY;
  wire CPLLLOCKDETCLK_INDELAY;
  wire CPLLLOCKEN_INDELAY;
  wire CPLLPD_INDELAY;
  wire CPLLRESET_INDELAY;
  wire DRPCLK_INDELAY;
  wire DRPEN_INDELAY;
  wire DRPWE_INDELAY;
  wire EYESCANMODE_INDELAY;
  wire EYESCANRESET_INDELAY;
  wire EYESCANTRIGGER_INDELAY;
  wire GTGREFCLK_INDELAY;
  wire GTNORTHREFCLK0_INDELAY;
  wire GTNORTHREFCLK1_INDELAY;
  wire GTREFCLK0_INDELAY;
  wire GTREFCLK1_INDELAY;
  wire GTRESETSEL_INDELAY;
  wire GTRXRESET_INDELAY;
  wire GTSOUTHREFCLK0_INDELAY;
  wire GTSOUTHREFCLK1_INDELAY;
  wire GTTXRESET_INDELAY;
  wire GTXRXN_INDELAY;
  wire GTXRXP_INDELAY;
  wire QPLLCLK_INDELAY;
  wire QPLLREFCLK_INDELAY;
  wire RESETOVRD_INDELAY;
  wire RX8B10BEN_INDELAY;
  wire RXBUFRESET_INDELAY;
  wire RXCDRFREQRESET_INDELAY;
  wire RXCDRHOLD_INDELAY;
  wire RXCDROVRDEN_INDELAY;
  wire RXCDRRESETRSV_INDELAY;
  wire RXCDRRESET_INDELAY;
  wire RXCHBONDEN_INDELAY;
  wire RXCHBONDMASTER_INDELAY;
  wire RXCHBONDSLAVE_INDELAY;
  wire RXCOMMADETEN_INDELAY;
  wire RXDDIEN_INDELAY;
  wire RXDFEAGCHOLD_INDELAY;
  wire RXDFEAGCOVRDEN_INDELAY;
  wire RXDFECM1EN_INDELAY;
  wire RXDFELFHOLD_INDELAY;
  wire RXDFELFOVRDEN_INDELAY;
  wire RXDFELPMRESET_INDELAY;
  wire RXDFETAP2HOLD_INDELAY;
  wire RXDFETAP2OVRDEN_INDELAY;
  wire RXDFETAP3HOLD_INDELAY;
  wire RXDFETAP3OVRDEN_INDELAY;
  wire RXDFETAP4HOLD_INDELAY;
  wire RXDFETAP4OVRDEN_INDELAY;
  wire RXDFETAP5HOLD_INDELAY;
  wire RXDFETAP5OVRDEN_INDELAY;
  wire RXDFEUTHOLD_INDELAY;
  wire RXDFEUTOVRDEN_INDELAY;
  wire RXDFEVPHOLD_INDELAY;
  wire RXDFEVPOVRDEN_INDELAY;
  wire RXDFEVSEN_INDELAY;
  wire RXDFEXYDEN_INDELAY;
  wire RXDFEXYDHOLD_INDELAY;
  wire RXDFEXYDOVRDEN_INDELAY;
  wire RXDLYBYPASS_INDELAY;
  wire RXDLYEN_INDELAY;
  wire RXDLYOVRDEN_INDELAY;
  wire RXDLYSRESET_INDELAY;
  wire RXGEARBOXSLIP_INDELAY;
  wire RXLPMEN_INDELAY;
  wire RXLPMHFHOLD_INDELAY;
  wire RXLPMHFOVRDEN_INDELAY;
  wire RXLPMLFHOLD_INDELAY;
  wire RXLPMLFKLOVRDEN_INDELAY;
  wire RXMCOMMAALIGNEN_INDELAY;
  wire RXOOBRESET_INDELAY;
  wire RXOSHOLD_INDELAY;
  wire RXOSOVRDEN_INDELAY;
  wire RXPCOMMAALIGNEN_INDELAY;
  wire RXPCSRESET_INDELAY;
  wire RXPHALIGNEN_INDELAY;
  wire RXPHALIGN_INDELAY;
  wire RXPHDLYPD_INDELAY;
  wire RXPHDLYRESET_INDELAY;
  wire RXPHOVRDEN_INDELAY;
  wire RXPMARESET_INDELAY;
  wire RXPOLARITY_INDELAY;
  wire RXPRBSCNTRESET_INDELAY;
  wire RXQPIEN_INDELAY;
  wire RXSLIDE_INDELAY;
  wire RXUSERRDY_INDELAY;
  wire RXUSRCLK2_INDELAY;
  wire RXUSRCLK_INDELAY;
  wire SETERRSTATUS_INDELAY;
  wire TX8B10BEN_INDELAY;
  wire TXCOMINIT_INDELAY;
  wire TXCOMSAS_INDELAY;
  wire TXCOMWAKE_INDELAY;
  wire TXDEEMPH_INDELAY;
  wire TXDETECTRX_INDELAY;
  wire TXDIFFPD_INDELAY;
  wire TXDLYBYPASS_INDELAY;
  wire TXDLYEN_INDELAY;
  wire TXDLYHOLD_INDELAY;
  wire TXDLYOVRDEN_INDELAY;
  wire TXDLYSRESET_INDELAY;
  wire TXDLYUPDOWN_INDELAY;
  wire TXELECIDLE_INDELAY;
  wire TXINHIBIT_INDELAY;
  wire TXPCSRESET_INDELAY;
  wire TXPDELECIDLEMODE_INDELAY;
  wire TXPHALIGNEN_INDELAY;
  wire TXPHALIGN_INDELAY;
  wire TXPHDLYPD_INDELAY;
  wire TXPHDLYRESET_INDELAY;
  wire TXPHDLYTSTCLK_INDELAY;
  wire TXPHINIT_INDELAY;
  wire TXPHOVRDEN_INDELAY;
  wire TXPISOPD_INDELAY;
  wire TXPMARESET_INDELAY;
  wire TXPOLARITY_INDELAY;
  wire TXPOSTCURSORINV_INDELAY;
  wire TXPRBSFORCEERR_INDELAY;
  wire TXPRECURSORINV_INDELAY;
  wire TXQPIBIASEN_INDELAY;
  wire TXQPISTRONGPDOWN_INDELAY;
  wire TXQPIWEAKPUP_INDELAY;
  wire TXSTARTSEQ_INDELAY;
  wire TXSWING_INDELAY;
  wire TXUSERRDY_INDELAY;
  wire TXUSRCLK2_INDELAY;
  wire TXUSRCLK_INDELAY;
  wire [15:0] DRPDI_INDELAY;
  wire [15:0] GTRSVD_INDELAY;
  wire [15:0] PCSRSVDIN_INDELAY;
  wire [19:0] TSTIN_INDELAY;
  wire [1:0] RXELECIDLEMODE_INDELAY;
  wire [1:0] RXMONITORSEL_INDELAY;
  wire [1:0] RXPD_INDELAY;
  wire [1:0] RXSYSCLKSEL_INDELAY;
  wire [1:0] TXPD_INDELAY;
  wire [1:0] TXSYSCLKSEL_INDELAY;
  wire [2:0] CPLLREFCLKSEL_INDELAY;
  wire [2:0] LOOPBACK_INDELAY;
  wire [2:0] RXCHBONDLEVEL_INDELAY;
  wire [2:0] RXOUTCLKSEL_INDELAY;
  wire [2:0] RXPRBSSEL_INDELAY;
  wire [2:0] RXRATE_INDELAY;
  wire [2:0] TXBUFDIFFCTRL_INDELAY;
  wire [2:0] TXHEADER_INDELAY;
  wire [2:0] TXMARGIN_INDELAY;
  wire [2:0] TXOUTCLKSEL_INDELAY;
  wire [2:0] TXPRBSSEL_INDELAY;
  wire [2:0] TXRATE_INDELAY;
  wire [3:0] CLKRSVD_INDELAY;
  wire [3:0] TXDIFFCTRL_INDELAY;
  wire [4:0] PCSRSVDIN2_INDELAY;
  wire [4:0] PMARSVDIN2_INDELAY;
  wire [4:0] PMARSVDIN_INDELAY;
  wire [4:0] RXCHBONDI_INDELAY;
  wire [4:0] TXPOSTCURSOR_INDELAY;
  wire [4:0] TXPRECURSOR_INDELAY;
  wire [63:0] TXDATA_INDELAY;
  wire [6:0] TXMAINCURSOR_INDELAY;
  wire [6:0] TXSEQUENCE_INDELAY;
  wire [7:0] TX8B10BBYPASS_INDELAY;
  wire [7:0] TXCHARDISPMODE_INDELAY;
  wire [7:0] TXCHARDISPVAL_INDELAY;
  wire [7:0] TXCHARISK_INDELAY;
  wire [8:0] DRPADDR_INDELAY;

  initial begin
    case (ALIGN_COMMA_DOUBLE)
      "FALSE" : ALIGN_COMMA_DOUBLE_BINARY = 1'b0;
      "TRUE" : ALIGN_COMMA_DOUBLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ALIGN_COMMA_DOUBLE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ALIGN_COMMA_DOUBLE);
        $finish;
      end
    endcase

    case (ALIGN_COMMA_WORD)
      1 : ALIGN_COMMA_WORD_BINARY = 3'b001;
      2 : ALIGN_COMMA_WORD_BINARY = 3'b010;
      4 : ALIGN_COMMA_WORD_BINARY = 3'b100;
      default : begin
        $display("Attribute Syntax Error : The Attribute ALIGN_COMMA_WORD on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 4.", ALIGN_COMMA_WORD, 1);
        $finish;
      end
    endcase

    case (ALIGN_MCOMMA_DET)
      "TRUE" : ALIGN_MCOMMA_DET_BINARY = 1'b1;
      "FALSE" : ALIGN_MCOMMA_DET_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute ALIGN_MCOMMA_DET on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", ALIGN_MCOMMA_DET);
        $finish;
      end
    endcase

    case (ALIGN_PCOMMA_DET)
      "TRUE" : ALIGN_PCOMMA_DET_BINARY = 1'b1;
      "FALSE" : ALIGN_PCOMMA_DET_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute ALIGN_PCOMMA_DET on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", ALIGN_PCOMMA_DET);
        $finish;
      end
    endcase

    case (CBCC_DATA_SOURCE_SEL)
      "DECODED" : CBCC_DATA_SOURCE_SEL_BINARY = 1'b1;
      "ENCODED" : CBCC_DATA_SOURCE_SEL_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CBCC_DATA_SOURCE_SEL on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are DECODED, or ENCODED.", CBCC_DATA_SOURCE_SEL);
        $finish;
      end
    endcase

    case (CHAN_BOND_KEEP_ALIGN)
      "FALSE" : CHAN_BOND_KEEP_ALIGN_BINARY = 1'b0;
      "TRUE" : CHAN_BOND_KEEP_ALIGN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute CHAN_BOND_KEEP_ALIGN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", CHAN_BOND_KEEP_ALIGN);
        $finish;
      end
    endcase

    case (CHAN_BOND_SEQ_2_USE)
      "FALSE" : CHAN_BOND_SEQ_2_USE_BINARY = 1'b0;
      "TRUE" : CHAN_BOND_SEQ_2_USE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_USE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", CHAN_BOND_SEQ_2_USE);
        $finish;
      end
    endcase

    case (CHAN_BOND_SEQ_LEN)
      1 : CHAN_BOND_SEQ_LEN_BINARY = 2'b00;
      2 : CHAN_BOND_SEQ_LEN_BINARY = 2'b01;
      3 : CHAN_BOND_SEQ_LEN_BINARY = 2'b10;
      4 : CHAN_BOND_SEQ_LEN_BINARY = 2'b11;
      default : begin
        $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_LEN on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 4.", CHAN_BOND_SEQ_LEN, 1);
        $finish;
      end
    endcase

    case (CLK_CORRECT_USE)
      "TRUE" : CLK_CORRECT_USE_BINARY = 1'b1;
      "FALSE" : CLK_CORRECT_USE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CLK_CORRECT_USE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", CLK_CORRECT_USE);
        $finish;
      end
    endcase

    case (CLK_COR_KEEP_IDLE)
      "FALSE" : CLK_COR_KEEP_IDLE_BINARY = 1'b0;
      "TRUE" : CLK_COR_KEEP_IDLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute CLK_COR_KEEP_IDLE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", CLK_COR_KEEP_IDLE);
        $finish;
      end
    endcase

    case (CLK_COR_PRECEDENCE)
      "TRUE" : CLK_COR_PRECEDENCE_BINARY = 1'b1;
      "FALSE" : CLK_COR_PRECEDENCE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CLK_COR_PRECEDENCE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", CLK_COR_PRECEDENCE);
        $finish;
      end
    endcase

    case (CLK_COR_SEQ_2_USE)
      "FALSE" : CLK_COR_SEQ_2_USE_BINARY = 1'b0;
      "TRUE" : CLK_COR_SEQ_2_USE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_USE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", CLK_COR_SEQ_2_USE);
        $finish;
      end
    endcase

    case (CLK_COR_SEQ_LEN)
      1 : CLK_COR_SEQ_LEN_BINARY = 2'b00;
      2 : CLK_COR_SEQ_LEN_BINARY = 2'b01;
      3 : CLK_COR_SEQ_LEN_BINARY = 2'b10;
      4 : CLK_COR_SEQ_LEN_BINARY = 2'b11;
      default : begin
        $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_LEN on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 4.", CLK_COR_SEQ_LEN, 1);
        $finish;
      end
    endcase

    case (CPLL_FBDIV)
      4 : CPLL_FBDIV_BINARY = 7'b0000010;
      1 : CPLL_FBDIV_BINARY = 7'b0010000;
      2 : CPLL_FBDIV_BINARY = 7'b0000000;
      3 : CPLL_FBDIV_BINARY = 7'b0000001;
      5 : CPLL_FBDIV_BINARY = 7'b0000011;
      6 : CPLL_FBDIV_BINARY = 7'b0000101;
      8 : CPLL_FBDIV_BINARY = 7'b0000110;
      10 : CPLL_FBDIV_BINARY = 7'b0000111;
      12 : CPLL_FBDIV_BINARY = 7'b0001101;
      16 : CPLL_FBDIV_BINARY = 7'b0001110;
      20 : CPLL_FBDIV_BINARY = 7'b0001111;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPLL_FBDIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 20.", CPLL_FBDIV, 4);
        $finish;
      end
    endcase

    case (CPLL_FBDIV_45)
      5 : CPLL_FBDIV_45_BINARY = 1'b1;
      4 : CPLL_FBDIV_45_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPLL_FBDIV_45 on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 4 to 5.", CPLL_FBDIV_45, 5);
        $finish;
      end
    endcase

    case (CPLL_REFCLK_DIV)
      1 : CPLL_REFCLK_DIV_BINARY = 5'b10000;
      2 : CPLL_REFCLK_DIV_BINARY = 5'b00000;
      3 : CPLL_REFCLK_DIV_BINARY = 5'b00001;
      4 : CPLL_REFCLK_DIV_BINARY = 5'b00010;
      5 : CPLL_REFCLK_DIV_BINARY = 5'b00011;
      6 : CPLL_REFCLK_DIV_BINARY = 5'b00101;
      8 : CPLL_REFCLK_DIV_BINARY = 5'b00110;
      10 : CPLL_REFCLK_DIV_BINARY = 5'b00111;
      12 : CPLL_REFCLK_DIV_BINARY = 5'b01101;
      16 : CPLL_REFCLK_DIV_BINARY = 5'b01110;
      20 : CPLL_REFCLK_DIV_BINARY = 5'b01111;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPLL_REFCLK_DIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 20.", CPLL_REFCLK_DIV, 1);
        $finish;
      end
    endcase

    case (CPLL_RXOUT_DIV)
      2 : CPLL_RXOUT_DIV_BINARY = 3'b001;
      1 : CPLL_RXOUT_DIV_BINARY = 3'b000;
      4 : CPLL_RXOUT_DIV_BINARY = 3'b010;
      8 : CPLL_RXOUT_DIV_BINARY = 3'b011;
      16 : CPLL_RXOUT_DIV_BINARY = 3'b100;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPLL_RXOUT_DIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 16.", CPLL_RXOUT_DIV, 2);
        $finish;
      end
    endcase

    case (CPLL_TXOUT_DIV)
      2 : CPLL_TXOUT_DIV_BINARY = 3'b001;
      1 : CPLL_TXOUT_DIV_BINARY = 3'b000;
      4 : CPLL_TXOUT_DIV_BINARY = 3'b010;
      8 : CPLL_TXOUT_DIV_BINARY = 3'b011;
      16 : CPLL_TXOUT_DIV_BINARY = 3'b100;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPLL_TXOUT_DIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 16.", CPLL_TXOUT_DIV, 2);
        $finish;
      end
    endcase

    case (DEC_MCOMMA_DETECT)
      "TRUE" : DEC_MCOMMA_DETECT_BINARY = 1'b1;
      "FALSE" : DEC_MCOMMA_DETECT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEC_MCOMMA_DETECT on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEC_MCOMMA_DETECT);
        $finish;
      end
    endcase

    case (DEC_PCOMMA_DETECT)
      "TRUE" : DEC_PCOMMA_DETECT_BINARY = 1'b1;
      "FALSE" : DEC_PCOMMA_DETECT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEC_PCOMMA_DETECT on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEC_PCOMMA_DETECT);
        $finish;
      end
    endcase

    case (DEC_VALID_COMMA_ONLY)
      "TRUE" : DEC_VALID_COMMA_ONLY_BINARY = 1'b1;
      "FALSE" : DEC_VALID_COMMA_ONLY_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEC_VALID_COMMA_ONLY on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEC_VALID_COMMA_ONLY);
        $finish;
      end
    endcase

    case (ES_ERRDET_EN)
      "FALSE" : ES_ERRDET_EN_BINARY = 1'b0;
      "TRUE" : ES_ERRDET_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ES_ERRDET_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ES_ERRDET_EN);
        $finish;
      end
    endcase

    case (ES_EYE_SCAN_EN)
      "FALSE" : ES_EYE_SCAN_EN_BINARY = 1'b0;
      "TRUE" : ES_EYE_SCAN_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ES_EYE_SCAN_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ES_EYE_SCAN_EN);
        $finish;
      end
    endcase

    case (FTS_LANE_DESKEW_EN)
      "FALSE" : FTS_LANE_DESKEW_EN_BINARY = 1'b0;
      "TRUE" : FTS_LANE_DESKEW_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute FTS_LANE_DESKEW_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", FTS_LANE_DESKEW_EN);
        $finish;
      end
    endcase

    case (PCS_PCIE_EN)
      "FALSE" : PCS_PCIE_EN_BINARY = 1'b0;
      "TRUE" : PCS_PCIE_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PCS_PCIE_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PCS_PCIE_EN);
        $finish;
      end
    endcase

    case (RXBUF_ADDR_MODE)
      "FULL" : RXBUF_ADDR_MODE_BINARY = 1'b0;
      "FAST" : RXBUF_ADDR_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_ADDR_MODE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FULL, or FAST.", RXBUF_ADDR_MODE);
        $finish;
      end
    endcase

    case (RXBUF_EN)
      "TRUE" : RXBUF_EN_BINARY = 1'b1;
      "FALSE" : RXBUF_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RXBUF_EN);
        $finish;
      end
    endcase

    case (RXBUF_RESET_ON_CB_CHANGE)
      "TRUE" : RXBUF_RESET_ON_CB_CHANGE_BINARY = 1'b1;
      "FALSE" : RXBUF_RESET_ON_CB_CHANGE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_RESET_ON_CB_CHANGE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RXBUF_RESET_ON_CB_CHANGE);
        $finish;
      end
    endcase

    case (RXBUF_RESET_ON_COMMAALIGN)
      "FALSE" : RXBUF_RESET_ON_COMMAALIGN_BINARY = 1'b0;
      "TRUE" : RXBUF_RESET_ON_COMMAALIGN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_RESET_ON_COMMAALIGN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", RXBUF_RESET_ON_COMMAALIGN);
        $finish;
      end
    endcase

    case (RXBUF_RESET_ON_EIDLE)
      "TRUE" : RXBUF_RESET_ON_EIDLE_BINARY = 1'b1;
      "FALSE" : RXBUF_RESET_ON_EIDLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_RESET_ON_EIDLE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RXBUF_RESET_ON_EIDLE);
        $finish;
      end
    endcase

    case (RXBUF_RESET_ON_RATE_CHANGE)
      "TRUE" : RXBUF_RESET_ON_RATE_CHANGE_BINARY = 1'b1;
      "FALSE" : RXBUF_RESET_ON_RATE_CHANGE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_RESET_ON_RATE_CHANGE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RXBUF_RESET_ON_RATE_CHANGE);
        $finish;
      end
    endcase

    case (RXBUF_THRESH_OVRD)
      "FALSE" : RXBUF_THRESH_OVRD_BINARY = 1'b0;
      "TRUE" : RXBUF_THRESH_OVRD_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXBUF_THRESH_OVRD on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", RXBUF_THRESH_OVRD);
        $finish;
      end
    endcase

    case (RXGEARBOX_EN)
      "FALSE" : RXGEARBOX_EN_BINARY = 1'b0;
      "TRUE" : RXGEARBOX_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXGEARBOX_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", RXGEARBOX_EN);
        $finish;
      end
    endcase

    case (RXSLIDE_MODE)
      "OFF" : RXSLIDE_MODE_BINARY = 2'b00;
      "AUTO" : RXSLIDE_MODE_BINARY = 2'b01;
      "PCS" : RXSLIDE_MODE_BINARY = 2'b10;
      "PMA" : RXSLIDE_MODE_BINARY = 2'b11;
      default : begin
        $display("Attribute Syntax Error : The Attribute RXSLIDE_MODE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are OFF, AUTO, PCS, or PMA.", RXSLIDE_MODE);
        $finish;
      end
    endcase

    case (RX_CLK25_DIV)
      7 : RX_CLK25_DIV_BINARY = 5'b00110;
      1 : RX_CLK25_DIV_BINARY = 5'b00000;
      2 : RX_CLK25_DIV_BINARY = 5'b00001;
      3 : RX_CLK25_DIV_BINARY = 5'b00010;
      4 : RX_CLK25_DIV_BINARY = 5'b00011;
      5 : RX_CLK25_DIV_BINARY = 5'b00100;
      6 : RX_CLK25_DIV_BINARY = 5'b00101;
      8 : RX_CLK25_DIV_BINARY = 5'b00111;
      9 : RX_CLK25_DIV_BINARY = 5'b01000;
      10 : RX_CLK25_DIV_BINARY = 5'b01001;
      11 : RX_CLK25_DIV_BINARY = 5'b01010;
      12 : RX_CLK25_DIV_BINARY = 5'b01011;
      13 : RX_CLK25_DIV_BINARY = 5'b01100;
      14 : RX_CLK25_DIV_BINARY = 5'b01101;
      15 : RX_CLK25_DIV_BINARY = 5'b01110;
      16 : RX_CLK25_DIV_BINARY = 5'b01111;
      17 : RX_CLK25_DIV_BINARY = 5'b10000;
      18 : RX_CLK25_DIV_BINARY = 5'b10001;
      19 : RX_CLK25_DIV_BINARY = 5'b10010;
      20 : RX_CLK25_DIV_BINARY = 5'b10011;
      21 : RX_CLK25_DIV_BINARY = 5'b10100;
      22 : RX_CLK25_DIV_BINARY = 5'b10101;
      23 : RX_CLK25_DIV_BINARY = 5'b10110;
      24 : RX_CLK25_DIV_BINARY = 5'b10111;
      25 : RX_CLK25_DIV_BINARY = 5'b11000;
      26 : RX_CLK25_DIV_BINARY = 5'b11001;
      27 : RX_CLK25_DIV_BINARY = 5'b11010;
      28 : RX_CLK25_DIV_BINARY = 5'b11011;
      29 : RX_CLK25_DIV_BINARY = 5'b11100;
      30 : RX_CLK25_DIV_BINARY = 5'b11101;
      31 : RX_CLK25_DIV_BINARY = 5'b11110;
      32 : RX_CLK25_DIV_BINARY = 5'b11111;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_CLK25_DIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 32.", RX_CLK25_DIV, 7);
        $finish;
      end
    endcase

    case (RX_DATA_WIDTH)
      20 : RX_DATA_WIDTH_BINARY = 3'b011;
      16 : RX_DATA_WIDTH_BINARY = 3'b010;
      32 : RX_DATA_WIDTH_BINARY = 3'b100;
      40 : RX_DATA_WIDTH_BINARY = 3'b101;
      64 : RX_DATA_WIDTH_BINARY = 3'b110;
      80 : RX_DATA_WIDTH_BINARY = 3'b111;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_DATA_WIDTH on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 16 to 80.", RX_DATA_WIDTH, 20);
        $finish;
      end
    endcase

    case (RX_DEFER_RESET_BUF_EN)
      "TRUE" : RX_DEFER_RESET_BUF_EN_BINARY = 1'b1;
      "FALSE" : RX_DEFER_RESET_BUF_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_DEFER_RESET_BUF_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RX_DEFER_RESET_BUF_EN);
        $finish;
      end
    endcase

    case (RX_DISPERR_SEQ_MATCH)
      "TRUE" : RX_DISPERR_SEQ_MATCH_BINARY = 1'b1;
      "FALSE" : RX_DISPERR_SEQ_MATCH_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_DISPERR_SEQ_MATCH on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", RX_DISPERR_SEQ_MATCH);
        $finish;
      end
    endcase

    case (RX_SIG_VALID_DLY)
      10 : RX_SIG_VALID_DLY_BINARY = 5'b01001;
      1 : RX_SIG_VALID_DLY_BINARY = 5'b00000;
      2 : RX_SIG_VALID_DLY_BINARY = 5'b00001;
      3 : RX_SIG_VALID_DLY_BINARY = 5'b00010;
      4 : RX_SIG_VALID_DLY_BINARY = 5'b00011;
      5 : RX_SIG_VALID_DLY_BINARY = 5'b00100;
      6 : RX_SIG_VALID_DLY_BINARY = 5'b00101;
      7 : RX_SIG_VALID_DLY_BINARY = 5'b00110;
      8 : RX_SIG_VALID_DLY_BINARY = 5'b00111;
      9 : RX_SIG_VALID_DLY_BINARY = 5'b01000;
      11 : RX_SIG_VALID_DLY_BINARY = 5'b01010;
      12 : RX_SIG_VALID_DLY_BINARY = 5'b01011;
      13 : RX_SIG_VALID_DLY_BINARY = 5'b01100;
      14 : RX_SIG_VALID_DLY_BINARY = 5'b01101;
      15 : RX_SIG_VALID_DLY_BINARY = 5'b01110;
      16 : RX_SIG_VALID_DLY_BINARY = 5'b01111;
      17 : RX_SIG_VALID_DLY_BINARY = 5'b10000;
      18 : RX_SIG_VALID_DLY_BINARY = 5'b10001;
      19 : RX_SIG_VALID_DLY_BINARY = 5'b10010;
      20 : RX_SIG_VALID_DLY_BINARY = 5'b10011;
      21 : RX_SIG_VALID_DLY_BINARY = 5'b10100;
      22 : RX_SIG_VALID_DLY_BINARY = 5'b10101;
      23 : RX_SIG_VALID_DLY_BINARY = 5'b10110;
      24 : RX_SIG_VALID_DLY_BINARY = 5'b10111;
      25 : RX_SIG_VALID_DLY_BINARY = 5'b11000;
      26 : RX_SIG_VALID_DLY_BINARY = 5'b11001;
      27 : RX_SIG_VALID_DLY_BINARY = 5'b11010;
      28 : RX_SIG_VALID_DLY_BINARY = 5'b11011;
      29 : RX_SIG_VALID_DLY_BINARY = 5'b11100;
      30 : RX_SIG_VALID_DLY_BINARY = 5'b11101;
      31 : RX_SIG_VALID_DLY_BINARY = 5'b11110;
      32 : RX_SIG_VALID_DLY_BINARY = 5'b11111;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_SIG_VALID_DLY on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 32.", RX_SIG_VALID_DLY, 10);
        $finish;
      end
    endcase

    case (RX_XCLK_SEL)
      "RXREC" : RX_XCLK_SEL_BINARY = 1'b0;
      "RXUSR" : RX_XCLK_SEL_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RX_XCLK_SEL on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are RXREC, or RXUSR.", RX_XCLK_SEL);
        $finish;
      end
    endcase

    case (SATA_CPLL_CFG)
      "VCO_3000MHZ" : SATA_CPLL_CFG_BINARY = 2'b00;
      "VCO_750MHZ" : SATA_CPLL_CFG_BINARY = 2'b10;
      "VCO_1500MHZ" : SATA_CPLL_CFG_BINARY = 2'b01;
      default : begin
        $display("Attribute Syntax Error : The Attribute SATA_CPLL_CFG on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are VCO_3000MHZ, VCO_750MHZ, or VCO_1500MHZ.", SATA_CPLL_CFG);
        $finish;
      end
    endcase

    case (SHOW_REALIGN_COMMA)
      "TRUE" : SHOW_REALIGN_COMMA_BINARY = 1'b1;
      "FALSE" : SHOW_REALIGN_COMMA_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SHOW_REALIGN_COMMA on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", SHOW_REALIGN_COMMA);
        $finish;
      end
    endcase

    case (SIM_RECEIVER_DETECT_PASS)
      "TRUE" : SIM_RECEIVER_DETECT_PASS_BINARY = 0;
      "FALSE" : SIM_RECEIVER_DETECT_PASS_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_RECEIVER_DETECT_PASS on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", SIM_RECEIVER_DETECT_PASS);
        $finish;
      end
    endcase

    case (SIM_RESET_SPEEDUP)
      "TRUE" : SIM_RESET_SPEEDUP_BINARY = 0;
      "FALSE" : SIM_RESET_SPEEDUP_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_RESET_SPEEDUP on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", SIM_RESET_SPEEDUP);
        $finish;
      end
    endcase

    case (SIM_TX_EIDLE_DRIVE_LEVEL)
      "X" : SIM_TX_EIDLE_DRIVE_LEVEL_BINARY = 0;
      "0" : SIM_TX_EIDLE_DRIVE_LEVEL_BINARY = 0;
      "1" : SIM_TX_EIDLE_DRIVE_LEVEL_BINARY = 0;
      "Z" : SIM_TX_EIDLE_DRIVE_LEVEL_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_TX_EIDLE_DRIVE_LEVEL on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are X, 0, 1, or Z.", SIM_TX_EIDLE_DRIVE_LEVEL);
        $finish;
      end
    endcase

    case (SIM_VERSION)
      "1.0" : SIM_VERSION_BINARY = 0;
      "2.0" : SIM_VERSION_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_VERSION on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are 1.0, or 2.0.", SIM_VERSION);
        $finish;
      end
    endcase

    case (TXBUF_EN)
      "TRUE" : TXBUF_EN_BINARY = 1'b1;
      "FALSE" : TXBUF_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TXBUF_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", TXBUF_EN);
        $finish;
      end
    endcase

    case (TXBUF_RESET_ON_RATE_CHANGE)
      "FALSE" : TXBUF_RESET_ON_RATE_CHANGE_BINARY = 1'b0;
      "TRUE" : TXBUF_RESET_ON_RATE_CHANGE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TXBUF_RESET_ON_RATE_CHANGE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TXBUF_RESET_ON_RATE_CHANGE);
        $finish;
      end
    endcase

    case (TXGEARBOX_EN)
      "FALSE" : TXGEARBOX_EN_BINARY = 1'b0;
      "TRUE" : TXGEARBOX_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TXGEARBOX_EN on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TXGEARBOX_EN);
        $finish;
      end
    endcase

    case (TX_CLK25_DIV)
      7 : TX_CLK25_DIV_BINARY = 5'b00110;
      1 : TX_CLK25_DIV_BINARY = 5'b00000;
      2 : TX_CLK25_DIV_BINARY = 5'b00001;
      3 : TX_CLK25_DIV_BINARY = 5'b00010;
      4 : TX_CLK25_DIV_BINARY = 5'b00011;
      5 : TX_CLK25_DIV_BINARY = 5'b00100;
      6 : TX_CLK25_DIV_BINARY = 5'b00101;
      8 : TX_CLK25_DIV_BINARY = 5'b00111;
      9 : TX_CLK25_DIV_BINARY = 5'b01000;
      10 : TX_CLK25_DIV_BINARY = 5'b01001;
      11 : TX_CLK25_DIV_BINARY = 5'b01010;
      12 : TX_CLK25_DIV_BINARY = 5'b01011;
      13 : TX_CLK25_DIV_BINARY = 5'b01100;
      14 : TX_CLK25_DIV_BINARY = 5'b01101;
      15 : TX_CLK25_DIV_BINARY = 5'b01110;
      16 : TX_CLK25_DIV_BINARY = 5'b01111;
      17 : TX_CLK25_DIV_BINARY = 5'b10000;
      18 : TX_CLK25_DIV_BINARY = 5'b10001;
      19 : TX_CLK25_DIV_BINARY = 5'b10010;
      20 : TX_CLK25_DIV_BINARY = 5'b10011;
      21 : TX_CLK25_DIV_BINARY = 5'b10100;
      22 : TX_CLK25_DIV_BINARY = 5'b10101;
      23 : TX_CLK25_DIV_BINARY = 5'b10110;
      24 : TX_CLK25_DIV_BINARY = 5'b10111;
      25 : TX_CLK25_DIV_BINARY = 5'b11000;
      26 : TX_CLK25_DIV_BINARY = 5'b11001;
      27 : TX_CLK25_DIV_BINARY = 5'b11010;
      28 : TX_CLK25_DIV_BINARY = 5'b11011;
      29 : TX_CLK25_DIV_BINARY = 5'b11100;
      30 : TX_CLK25_DIV_BINARY = 5'b11101;
      31 : TX_CLK25_DIV_BINARY = 5'b11110;
      32 : TX_CLK25_DIV_BINARY = 5'b11111;
      default : begin
        $display("Attribute Syntax Error : The Attribute TX_CLK25_DIV on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 1 to 32.", TX_CLK25_DIV, 7);
        $finish;
      end
    endcase

    case (TX_DATA_WIDTH)
      20 : TX_DATA_WIDTH_BINARY = 3'b011;
      16 : TX_DATA_WIDTH_BINARY = 3'b010;
      32 : TX_DATA_WIDTH_BINARY = 3'b100;
      40 : TX_DATA_WIDTH_BINARY = 3'b101;
      64 : TX_DATA_WIDTH_BINARY = 3'b110;
      80 : TX_DATA_WIDTH_BINARY = 3'b111;
      default : begin
        $display("Attribute Syntax Error : The Attribute TX_DATA_WIDTH on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are 16 to 80.", TX_DATA_WIDTH, 20);
        $finish;
      end
    endcase

    case (TX_DRIVE_MODE)
      "DIRECT" : TX_DRIVE_MODE_BINARY = 5'b00000;
      "PIPE" : TX_DRIVE_MODE_BINARY = 5'b00001;
      "PIPEGEN3" : TX_DRIVE_MODE_BINARY = 5'b00010;
      default : begin
        $display("Attribute Syntax Error : The Attribute TX_DRIVE_MODE on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are DIRECT, PIPE, or PIPEGEN3.", TX_DRIVE_MODE);
        $finish;
      end
    endcase

    case (TX_LOOPBACK_DRIVE_HIZ)
      "FALSE" : TX_LOOPBACK_DRIVE_HIZ_BINARY = 1'b0;
      "TRUE" : TX_LOOPBACK_DRIVE_HIZ_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TX_LOOPBACK_DRIVE_HIZ on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TX_LOOPBACK_DRIVE_HIZ);
        $finish;
      end
    endcase

    case (TX_XCLK_SEL)
      "TXUSR" : TX_XCLK_SEL_BINARY = 1'b1;
      "TXOUT" : TX_XCLK_SEL_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TX_XCLK_SEL on X_GTXE2_CHANNEL instance %m is set to %s.  Legal values for this attribute are TXUSR, or TXOUT.", TX_XCLK_SEL);
        $finish;
      end
    endcase

    if ((ALIGN_COMMA_ENABLE >= 10'b0000000000) && (ALIGN_COMMA_ENABLE <= 10'b1111111111))
      ALIGN_COMMA_ENABLE_BINARY = ALIGN_COMMA_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute ALIGN_COMMA_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", ALIGN_COMMA_ENABLE);
      $finish;
    end

    if ((ALIGN_MCOMMA_VALUE >= 10'b0000000000) && (ALIGN_MCOMMA_VALUE <= 10'b1111111111))
      ALIGN_MCOMMA_VALUE_BINARY = ALIGN_MCOMMA_VALUE;
    else begin
      $display("Attribute Syntax Error : The Attribute ALIGN_MCOMMA_VALUE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", ALIGN_MCOMMA_VALUE);
      $finish;
    end

    if ((ALIGN_PCOMMA_VALUE >= 10'b0000000000) && (ALIGN_PCOMMA_VALUE <= 10'b1111111111))
      ALIGN_PCOMMA_VALUE_BINARY = ALIGN_PCOMMA_VALUE;
    else begin
      $display("Attribute Syntax Error : The Attribute ALIGN_PCOMMA_VALUE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", ALIGN_PCOMMA_VALUE);
      $finish;
    end

    if ((CHAN_BOND_MAX_SKEW >= 1) && (CHAN_BOND_MAX_SKEW <= 14))
      CHAN_BOND_MAX_SKEW_BINARY = CHAN_BOND_MAX_SKEW;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_MAX_SKEW on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 14.", CHAN_BOND_MAX_SKEW);
      $finish;
    end

    if ((CHAN_BOND_SEQ_1_1 >= 10'b0000000000) && (CHAN_BOND_SEQ_1_1 <= 10'b1111111111))
      CHAN_BOND_SEQ_1_1_BINARY = CHAN_BOND_SEQ_1_1;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_1_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_1_1);
      $finish;
    end

    if ((CHAN_BOND_SEQ_1_2 >= 10'b0000000000) && (CHAN_BOND_SEQ_1_2 <= 10'b1111111111))
      CHAN_BOND_SEQ_1_2_BINARY = CHAN_BOND_SEQ_1_2;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_1_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_1_2);
      $finish;
    end

    if ((CHAN_BOND_SEQ_1_3 >= 10'b0000000000) && (CHAN_BOND_SEQ_1_3 <= 10'b1111111111))
      CHAN_BOND_SEQ_1_3_BINARY = CHAN_BOND_SEQ_1_3;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_1_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_1_3);
      $finish;
    end

    if ((CHAN_BOND_SEQ_1_4 >= 10'b0000000000) && (CHAN_BOND_SEQ_1_4 <= 10'b1111111111))
      CHAN_BOND_SEQ_1_4_BINARY = CHAN_BOND_SEQ_1_4;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_1_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_1_4);
      $finish;
    end

    if ((CHAN_BOND_SEQ_1_ENABLE >= 4'b0000) && (CHAN_BOND_SEQ_1_ENABLE <= 4'b1111))
      CHAN_BOND_SEQ_1_ENABLE_BINARY = CHAN_BOND_SEQ_1_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_1_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", CHAN_BOND_SEQ_1_ENABLE);
      $finish;
    end

    if ((CHAN_BOND_SEQ_2_1 >= 10'b0000000000) && (CHAN_BOND_SEQ_2_1 <= 10'b1111111111))
      CHAN_BOND_SEQ_2_1_BINARY = CHAN_BOND_SEQ_2_1;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_2_1);
      $finish;
    end

    if ((CHAN_BOND_SEQ_2_2 >= 10'b0000000000) && (CHAN_BOND_SEQ_2_2 <= 10'b1111111111))
      CHAN_BOND_SEQ_2_2_BINARY = CHAN_BOND_SEQ_2_2;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_2_2);
      $finish;
    end

    if ((CHAN_BOND_SEQ_2_3 >= 10'b0000000000) && (CHAN_BOND_SEQ_2_3 <= 10'b1111111111))
      CHAN_BOND_SEQ_2_3_BINARY = CHAN_BOND_SEQ_2_3;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_2_3);
      $finish;
    end

    if ((CHAN_BOND_SEQ_2_4 >= 10'b0000000000) && (CHAN_BOND_SEQ_2_4 <= 10'b1111111111))
      CHAN_BOND_SEQ_2_4_BINARY = CHAN_BOND_SEQ_2_4;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CHAN_BOND_SEQ_2_4);
      $finish;
    end

    if ((CHAN_BOND_SEQ_2_ENABLE >= 4'b0000) && (CHAN_BOND_SEQ_2_ENABLE <= 4'b1111))
      CHAN_BOND_SEQ_2_ENABLE_BINARY = CHAN_BOND_SEQ_2_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute CHAN_BOND_SEQ_2_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", CHAN_BOND_SEQ_2_ENABLE);
      $finish;
    end

    if ((CLK_COR_MAX_LAT >= 3) && (CLK_COR_MAX_LAT <= 60))
      CLK_COR_MAX_LAT_BINARY = CLK_COR_MAX_LAT;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_MAX_LAT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  3 to 60.", CLK_COR_MAX_LAT);
      $finish;
    end

    if ((CLK_COR_MIN_LAT >= 3) && (CLK_COR_MIN_LAT <= 60))
      CLK_COR_MIN_LAT_BINARY = CLK_COR_MIN_LAT;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_MIN_LAT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  3 to 60.", CLK_COR_MIN_LAT);
      $finish;
    end

    if ((CLK_COR_REPEAT_WAIT >= 0) && (CLK_COR_REPEAT_WAIT <= 31))
      CLK_COR_REPEAT_WAIT_BINARY = CLK_COR_REPEAT_WAIT;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_REPEAT_WAIT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 31.", CLK_COR_REPEAT_WAIT);
      $finish;
    end

    if ((CLK_COR_SEQ_1_1 >= 10'b0000000000) && (CLK_COR_SEQ_1_1 <= 10'b1111111111))
      CLK_COR_SEQ_1_1_BINARY = CLK_COR_SEQ_1_1;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_1_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_1_1);
      $finish;
    end

    if ((CLK_COR_SEQ_1_2 >= 10'b0000000000) && (CLK_COR_SEQ_1_2 <= 10'b1111111111))
      CLK_COR_SEQ_1_2_BINARY = CLK_COR_SEQ_1_2;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_1_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_1_2);
      $finish;
    end

    if ((CLK_COR_SEQ_1_3 >= 10'b0000000000) && (CLK_COR_SEQ_1_3 <= 10'b1111111111))
      CLK_COR_SEQ_1_3_BINARY = CLK_COR_SEQ_1_3;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_1_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_1_3);
      $finish;
    end

    if ((CLK_COR_SEQ_1_4 >= 10'b0000000000) && (CLK_COR_SEQ_1_4 <= 10'b1111111111))
      CLK_COR_SEQ_1_4_BINARY = CLK_COR_SEQ_1_4;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_1_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_1_4);
      $finish;
    end

    if ((CLK_COR_SEQ_1_ENABLE >= 4'b0000) && (CLK_COR_SEQ_1_ENABLE <= 4'b1111))
      CLK_COR_SEQ_1_ENABLE_BINARY = CLK_COR_SEQ_1_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_1_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", CLK_COR_SEQ_1_ENABLE);
      $finish;
    end

    if ((CLK_COR_SEQ_2_1 >= 10'b0000000000) && (CLK_COR_SEQ_2_1 <= 10'b1111111111))
      CLK_COR_SEQ_2_1_BINARY = CLK_COR_SEQ_2_1;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_2_1);
      $finish;
    end

    if ((CLK_COR_SEQ_2_2 >= 10'b0000000000) && (CLK_COR_SEQ_2_2 <= 10'b1111111111))
      CLK_COR_SEQ_2_2_BINARY = CLK_COR_SEQ_2_2;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_2_2);
      $finish;
    end

    if ((CLK_COR_SEQ_2_3 >= 10'b0000000000) && (CLK_COR_SEQ_2_3 <= 10'b1111111111))
      CLK_COR_SEQ_2_3_BINARY = CLK_COR_SEQ_2_3;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_2_3);
      $finish;
    end

    if ((CLK_COR_SEQ_2_4 >= 10'b0000000000) && (CLK_COR_SEQ_2_4 <= 10'b1111111111))
      CLK_COR_SEQ_2_4_BINARY = CLK_COR_SEQ_2_4;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", CLK_COR_SEQ_2_4);
      $finish;
    end

    if ((CLK_COR_SEQ_2_ENABLE >= 4'b0000) && (CLK_COR_SEQ_2_ENABLE <= 4'b1111))
      CLK_COR_SEQ_2_ENABLE_BINARY = CLK_COR_SEQ_2_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute CLK_COR_SEQ_2_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", CLK_COR_SEQ_2_ENABLE);
      $finish;
    end

    if ((ES_CONTROL >= 6'b000000) && (ES_CONTROL <= 6'b111111))
      ES_CONTROL_BINARY = ES_CONTROL;
    else begin
      $display("Attribute Syntax Error : The Attribute ES_CONTROL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 6'b000000 to 6'b111111.", ES_CONTROL);
      $finish;
    end

    if ((ES_PMA_CFG >= 10'b0000000000) && (ES_PMA_CFG <= 10'b1111111111))
      ES_PMA_CFG_BINARY = ES_PMA_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute ES_PMA_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 10'b0000000000 to 10'b1111111111.", ES_PMA_CFG);
      $finish;
    end

    if ((ES_PRESCALE >= 5'b00000) && (ES_PRESCALE <= 5'b11111))
      ES_PRESCALE_BINARY = ES_PRESCALE;
    else begin
      $display("Attribute Syntax Error : The Attribute ES_PRESCALE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", ES_PRESCALE);
      $finish;
    end

    if ((ES_VERT_OFFSET >= 9'b000000000) && (ES_VERT_OFFSET <= 9'b111111111))
      ES_VERT_OFFSET_BINARY = ES_VERT_OFFSET;
    else begin
      $display("Attribute Syntax Error : The Attribute ES_VERT_OFFSET on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 9'b000000000 to 9'b111111111.", ES_VERT_OFFSET);
      $finish;
    end

    if ((FTS_DESKEW_SEQ_ENABLE >= 4'b0000) && (FTS_DESKEW_SEQ_ENABLE <= 4'b1111))
      FTS_DESKEW_SEQ_ENABLE_BINARY = FTS_DESKEW_SEQ_ENABLE;
    else begin
      $display("Attribute Syntax Error : The Attribute FTS_DESKEW_SEQ_ENABLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", FTS_DESKEW_SEQ_ENABLE);
      $finish;
    end

    if ((FTS_LANE_DESKEW_CFG >= 4'b0000) && (FTS_LANE_DESKEW_CFG <= 4'b1111))
      FTS_LANE_DESKEW_CFG_BINARY = FTS_LANE_DESKEW_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute FTS_LANE_DESKEW_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", FTS_LANE_DESKEW_CFG);
      $finish;
    end

    if ((GEARBOX_MODE >= 3'b000) && (GEARBOX_MODE <= 3'b111))
      GEARBOX_MODE_BINARY = GEARBOX_MODE;
    else begin
      $display("Attribute Syntax Error : The Attribute GEARBOX_MODE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", GEARBOX_MODE);
      $finish;
    end

    if ((OUTREFCLK_SEL_INV >= 2'b00) && (OUTREFCLK_SEL_INV <= 2'b11))
      OUTREFCLK_SEL_INV_BINARY = OUTREFCLK_SEL_INV;
    else begin
      $display("Attribute Syntax Error : The Attribute OUTREFCLK_SEL_INV on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 2'b00 to 2'b11.", OUTREFCLK_SEL_INV);
      $finish;
    end

    if ((PMA_RSV3 >= 2'b00) && (PMA_RSV3 <= 2'b11))
      PMA_RSV3_BINARY = PMA_RSV3;
    else begin
      $display("Attribute Syntax Error : The Attribute PMA_RSV3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 2'b00 to 2'b11.", PMA_RSV3);
      $finish;
    end

    if ((RXBUFRESET_TIME >= 5'b00000) && (RXBUFRESET_TIME <= 5'b11111))
      RXBUFRESET_TIME_BINARY = RXBUFRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXBUFRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXBUFRESET_TIME);
      $finish;
    end

    if ((RXBUF_EIDLE_HI_CNT >= 4'b0000) && (RXBUF_EIDLE_HI_CNT <= 4'b1111))
      RXBUF_EIDLE_HI_CNT_BINARY = RXBUF_EIDLE_HI_CNT;
    else begin
      $display("Attribute Syntax Error : The Attribute RXBUF_EIDLE_HI_CNT on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", RXBUF_EIDLE_HI_CNT);
      $finish;
    end

    if ((RXBUF_EIDLE_LO_CNT >= 4'b0000) && (RXBUF_EIDLE_LO_CNT <= 4'b1111))
      RXBUF_EIDLE_LO_CNT_BINARY = RXBUF_EIDLE_LO_CNT;
    else begin
      $display("Attribute Syntax Error : The Attribute RXBUF_EIDLE_LO_CNT on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", RXBUF_EIDLE_LO_CNT);
      $finish;
    end

    if ((RXBUF_THRESH_OVFLW >= 0) && (RXBUF_THRESH_OVFLW <= 63))
      RXBUF_THRESH_OVFLW_BINARY = RXBUF_THRESH_OVFLW;
    else begin
      $display("Attribute Syntax Error : The Attribute RXBUF_THRESH_OVFLW on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 63.", RXBUF_THRESH_OVFLW);
      $finish;
    end

    if ((RXBUF_THRESH_UNDFLW >= 0) && (RXBUF_THRESH_UNDFLW <= 63))
      RXBUF_THRESH_UNDFLW_BINARY = RXBUF_THRESH_UNDFLW;
    else begin
      $display("Attribute Syntax Error : The Attribute RXBUF_THRESH_UNDFLW on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 63.", RXBUF_THRESH_UNDFLW);
      $finish;
    end

    if ((RXCDRFREQRESET_TIME >= 5'b00000) && (RXCDRFREQRESET_TIME <= 5'b11111))
      RXCDRFREQRESET_TIME_BINARY = RXCDRFREQRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDRFREQRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXCDRFREQRESET_TIME);
      $finish;
    end

    if ((RXCDRPHRESET_TIME >= 5'b00000) && (RXCDRPHRESET_TIME <= 5'b11111))
      RXCDRPHRESET_TIME_BINARY = RXCDRPHRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDRPHRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXCDRPHRESET_TIME);
      $finish;
    end

    if ((RXCDR_FR_RESET_ON_EIDLE >= 1'b0) && (RXCDR_FR_RESET_ON_EIDLE <= 1'b1))
      RXCDR_FR_RESET_ON_EIDLE_BINARY = RXCDR_FR_RESET_ON_EIDLE;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDR_FR_RESET_ON_EIDLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RXCDR_FR_RESET_ON_EIDLE);
      $finish;
    end

    if ((RXCDR_HOLD_DURING_EIDLE >= 1'b0) && (RXCDR_HOLD_DURING_EIDLE <= 1'b1))
      RXCDR_HOLD_DURING_EIDLE_BINARY = RXCDR_HOLD_DURING_EIDLE;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDR_HOLD_DURING_EIDLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RXCDR_HOLD_DURING_EIDLE);
      $finish;
    end

    if ((RXCDR_LOCK_CFG >= 6'b000000) && (RXCDR_LOCK_CFG <= 6'b111111))
      RXCDR_LOCK_CFG_BINARY = RXCDR_LOCK_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDR_LOCK_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 6'b000000 to 6'b111111.", RXCDR_LOCK_CFG);
      $finish;
    end

    if ((RXCDR_PH_RESET_ON_EIDLE >= 1'b0) && (RXCDR_PH_RESET_ON_EIDLE <= 1'b1))
      RXCDR_PH_RESET_ON_EIDLE_BINARY = RXCDR_PH_RESET_ON_EIDLE;
    else begin
      $display("Attribute Syntax Error : The Attribute RXCDR_PH_RESET_ON_EIDLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RXCDR_PH_RESET_ON_EIDLE);
      $finish;
    end

    if ((RXDFELPMRESET_TIME >= 7'b0000000) && (RXDFELPMRESET_TIME <= 7'b1111111))
      RXDFELPMRESET_TIME_BINARY = RXDFELPMRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXDFELPMRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", RXDFELPMRESET_TIME);
      $finish;
    end

    if ((RXISCANRESET_TIME >= 5'b00000) && (RXISCANRESET_TIME <= 5'b11111))
      RXISCANRESET_TIME_BINARY = RXISCANRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXISCANRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXISCANRESET_TIME);
      $finish;
    end

    if ((RXLPM_HF_CFG >= 14'b00000000000000) && (RXLPM_HF_CFG <= 14'b11111111111111))
      RXLPM_HF_CFG_BINARY = RXLPM_HF_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RXLPM_HF_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 14'b00000000000000 to 14'b11111111111111.", RXLPM_HF_CFG);
      $finish;
    end

    if ((RXLPM_LF_CFG >= 14'b00000000000000) && (RXLPM_LF_CFG <= 14'b11111111111111))
      RXLPM_LF_CFG_BINARY = RXLPM_LF_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RXLPM_LF_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 14'b00000000000000 to 14'b11111111111111.", RXLPM_LF_CFG);
      $finish;
    end

    if ((RXOOB_CFG >= 7'b0000000) && (RXOOB_CFG <= 7'b1111111))
      RXOOB_CFG_BINARY = RXOOB_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RXOOB_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", RXOOB_CFG);
      $finish;
    end

    if ((RXPCSRESET_TIME >= 5'b00000) && (RXPCSRESET_TIME <= 5'b11111))
      RXPCSRESET_TIME_BINARY = RXPCSRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXPCSRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXPCSRESET_TIME);
      $finish;
    end

    if ((RXPH_MONITOR_SEL >= 5'b00000) && (RXPH_MONITOR_SEL <= 5'b11111))
      RXPH_MONITOR_SEL_BINARY = RXPH_MONITOR_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute RXPH_MONITOR_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXPH_MONITOR_SEL);
      $finish;
    end

    if ((RXPMARESET_TIME >= 5'b00000) && (RXPMARESET_TIME <= 5'b11111))
      RXPMARESET_TIME_BINARY = RXPMARESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute RXPMARESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", RXPMARESET_TIME);
      $finish;
    end

    if ((RXPRBS_ERR_LOOPBACK >= 1'b0) && (RXPRBS_ERR_LOOPBACK <= 1'b1))
      RXPRBS_ERR_LOOPBACK_BINARY = RXPRBS_ERR_LOOPBACK;
    else begin
      $display("Attribute Syntax Error : The Attribute RXPRBS_ERR_LOOPBACK on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RXPRBS_ERR_LOOPBACK);
      $finish;
    end

    if ((RXSLIDE_AUTO_WAIT >= 0) && (RXSLIDE_AUTO_WAIT <= 15))
      RXSLIDE_AUTO_WAIT_BINARY = RXSLIDE_AUTO_WAIT;
    else begin
      $display("Attribute Syntax Error : The Attribute RXSLIDE_AUTO_WAIT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 15.", RXSLIDE_AUTO_WAIT);
      $finish;
    end

    if ((RX_BIAS_CFG >= 12'b000000000000) && (RX_BIAS_CFG <= 12'b111111111111))
      RX_BIAS_CFG_BINARY = RX_BIAS_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_BIAS_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 12'b000000000000 to 12'b111111111111.", RX_BIAS_CFG);
      $finish;
    end

    if ((RX_BUFFER_CFG >= 6'b000000) && (RX_BUFFER_CFG <= 6'b111111))
      RX_BUFFER_CFG_BINARY = RX_BUFFER_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_BUFFER_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 6'b000000 to 6'b111111.", RX_BUFFER_CFG);
      $finish;
    end

    if ((RX_CLKMUX_PD >= 1'b0) && (RX_CLKMUX_PD <= 1'b1))
      RX_CLKMUX_PD_BINARY = RX_CLKMUX_PD;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_CLKMUX_PD on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RX_CLKMUX_PD);
      $finish;
    end

    if ((RX_CM_SEL >= 2'b00) && (RX_CM_SEL <= 2'b11))
      RX_CM_SEL_BINARY = RX_CM_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_CM_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 2'b00 to 2'b11.", RX_CM_SEL);
      $finish;
    end

    if ((RX_CM_TRIM >= 3'b000) && (RX_CM_TRIM <= 3'b111))
      RX_CM_TRIM_BINARY = RX_CM_TRIM;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_CM_TRIM on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", RX_CM_TRIM);
      $finish;
    end

    if ((RX_DDI_SEL >= 6'b000000) && (RX_DDI_SEL <= 6'b111111))
      RX_DDI_SEL_BINARY = RX_DDI_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DDI_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 6'b000000 to 6'b111111.", RX_DDI_SEL);
      $finish;
    end

    if ((RX_DEBUG_CFG >= 12'b000000000000) && (RX_DEBUG_CFG <= 12'b111111111111))
      RX_DEBUG_CFG_BINARY = RX_DEBUG_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DEBUG_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 12'b000000000000 to 12'b111111111111.", RX_DEBUG_CFG);
      $finish;
    end

    if ((RX_DFE_H2_CFG >= 12'b000000000000) && (RX_DFE_H2_CFG <= 12'b111111111111))
      RX_DFE_H2_CFG_BINARY = RX_DFE_H2_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_H2_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 12'b000000000000 to 12'b111111111111.", RX_DFE_H2_CFG);
      $finish;
    end

    if ((RX_DFE_H3_CFG >= 12'b000000000000) && (RX_DFE_H3_CFG <= 12'b111111111111))
      RX_DFE_H3_CFG_BINARY = RX_DFE_H3_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_H3_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 12'b000000000000 to 12'b111111111111.", RX_DFE_H3_CFG);
      $finish;
    end

    if ((RX_DFE_H4_CFG >= 11'b00000000000) && (RX_DFE_H4_CFG <= 11'b11111111111))
      RX_DFE_H4_CFG_BINARY = RX_DFE_H4_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_H4_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 11'b00000000000 to 11'b11111111111.", RX_DFE_H4_CFG);
      $finish;
    end

    if ((RX_DFE_H5_CFG >= 11'b00000000000) && (RX_DFE_H5_CFG <= 11'b11111111111))
      RX_DFE_H5_CFG_BINARY = RX_DFE_H5_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_H5_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 11'b00000000000 to 11'b11111111111.", RX_DFE_H5_CFG);
      $finish;
    end

    if ((RX_DFE_KL_CFG >= 13'b0000000000000) && (RX_DFE_KL_CFG <= 13'b1111111111111))
      RX_DFE_KL_CFG_BINARY = RX_DFE_KL_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_KL_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 13'b0000000000000 to 13'b1111111111111.", RX_DFE_KL_CFG);
      $finish;
    end

    if ((RX_DFE_LPM_HOLD_DURING_EIDLE >= 1'b0) && (RX_DFE_LPM_HOLD_DURING_EIDLE <= 1'b1))
      RX_DFE_LPM_HOLD_DURING_EIDLE_BINARY = RX_DFE_LPM_HOLD_DURING_EIDLE;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_LPM_HOLD_DURING_EIDLE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", RX_DFE_LPM_HOLD_DURING_EIDLE);
      $finish;
    end

    if ((RX_DFE_UT_CFG >= 17'b00000000000000000) && (RX_DFE_UT_CFG <= 17'b11111111111111111))
      RX_DFE_UT_CFG_BINARY = RX_DFE_UT_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_UT_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 17'b00000000000000000 to 17'b11111111111111111.", RX_DFE_UT_CFG);
      $finish;
    end

    if ((RX_DFE_VP_CFG >= 17'b00000000000000000) && (RX_DFE_VP_CFG <= 17'b11111111111111111))
      RX_DFE_VP_CFG_BINARY = RX_DFE_VP_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_VP_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 17'b00000000000000000 to 17'b11111111111111111.", RX_DFE_VP_CFG);
      $finish;
    end

    if ((RX_DFE_XYD_CFG >= 13'b0000000000000) && (RX_DFE_XYD_CFG <= 13'b1111111111111))
      RX_DFE_XYD_CFG_BINARY = RX_DFE_XYD_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_DFE_XYD_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 13'b0000000000000 to 13'b1111111111111.", RX_DFE_XYD_CFG);
      $finish;
    end

    if ((RX_INT_DATAWIDTH >= 0) && (RX_INT_DATAWIDTH <= 1))
      RX_INT_DATAWIDTH_BINARY = RX_INT_DATAWIDTH;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_INT_DATAWIDTH on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 1.", RX_INT_DATAWIDTH);
      $finish;
    end

    if ((RX_OS_CFG >= 13'b0000000000000) && (RX_OS_CFG <= 13'b1111111111111))
      RX_OS_CFG_BINARY = RX_OS_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute RX_OS_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 13'b0000000000000 to 13'b1111111111111.", RX_OS_CFG);
      $finish;
    end

    if ((SAS_MAX_COM >= 1) && (SAS_MAX_COM <= 127))
      SAS_MAX_COM_BINARY = SAS_MAX_COM;
    else begin
      $display("Attribute Syntax Error : The Attribute SAS_MAX_COM on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 127.", SAS_MAX_COM);
      $finish;
    end

    if ((SAS_MIN_COM >= 1) && (SAS_MIN_COM <= 63))
      SAS_MIN_COM_BINARY = SAS_MIN_COM;
    else begin
      $display("Attribute Syntax Error : The Attribute SAS_MIN_COM on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SAS_MIN_COM);
      $finish;
    end

    if ((SATA_BURST_SEQ_LEN >= 4'b0000) && (SATA_BURST_SEQ_LEN <= 4'b1111))
      SATA_BURST_SEQ_LEN_BINARY = SATA_BURST_SEQ_LEN;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_BURST_SEQ_LEN on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 4'b0000 to 4'b1111.", SATA_BURST_SEQ_LEN);
      $finish;
    end

    if ((SATA_BURST_VAL >= 3'b000) && (SATA_BURST_VAL <= 3'b111))
      SATA_BURST_VAL_BINARY = SATA_BURST_VAL;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_BURST_VAL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", SATA_BURST_VAL);
      $finish;
    end

    if ((SATA_EIDLE_VAL >= 3'b000) && (SATA_EIDLE_VAL <= 3'b111))
      SATA_EIDLE_VAL_BINARY = SATA_EIDLE_VAL;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_EIDLE_VAL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", SATA_EIDLE_VAL);
      $finish;
    end

    if ((SATA_MAX_BURST >= 1) && (SATA_MAX_BURST <= 63))
      SATA_MAX_BURST_BINARY = SATA_MAX_BURST;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MAX_BURST on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SATA_MAX_BURST);
      $finish;
    end

    if ((SATA_MAX_INIT >= 1) && (SATA_MAX_INIT <= 63))
      SATA_MAX_INIT_BINARY = SATA_MAX_INIT;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MAX_INIT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SATA_MAX_INIT);
      $finish;
    end

    if ((SATA_MAX_WAKE >= 1) && (SATA_MAX_WAKE <= 63))
      SATA_MAX_WAKE_BINARY = SATA_MAX_WAKE;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MAX_WAKE on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SATA_MAX_WAKE);
      $finish;
    end

    if ((SATA_MIN_BURST >= 1) && (SATA_MIN_BURST <= 61))
      SATA_MIN_BURST_BINARY = SATA_MIN_BURST;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MIN_BURST on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 61.", SATA_MIN_BURST);
      $finish;
    end

    if ((SATA_MIN_INIT >= 1) && (SATA_MIN_INIT <= 63))
      SATA_MIN_INIT_BINARY = SATA_MIN_INIT;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MIN_INIT on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SATA_MIN_INIT);
      $finish;
    end

    if ((SATA_MIN_WAKE >= 1) && (SATA_MIN_WAKE <= 63))
      SATA_MIN_WAKE_BINARY = SATA_MIN_WAKE;
    else begin
      $display("Attribute Syntax Error : The Attribute SATA_MIN_WAKE on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  1 to 63.", SATA_MIN_WAKE);
      $finish;
    end

    if ((SIM_CPLLREFCLK_SEL >= 3'b0) && (SIM_CPLLREFCLK_SEL <= 3'b111))
      SIM_CPLLREFCLK_SEL_BINARY = SIM_CPLLREFCLK_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute SIM_CPLLREFCLK_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b0 to 3'b111.", SIM_CPLLREFCLK_SEL);
      $finish;
    end

    if ((TERM_RCAL_CFG >= 5'b00000) && (TERM_RCAL_CFG <= 5'b11111))
      TERM_RCAL_CFG_BINARY = TERM_RCAL_CFG;
    else begin
      $display("Attribute Syntax Error : The Attribute TERM_RCAL_CFG on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TERM_RCAL_CFG);
      $finish;
    end

    if ((TERM_RCAL_OVRD >= 1'b0) && (TERM_RCAL_OVRD <= 1'b1))
      TERM_RCAL_OVRD_BINARY = TERM_RCAL_OVRD;
    else begin
      $display("Attribute Syntax Error : The Attribute TERM_RCAL_OVRD on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", TERM_RCAL_OVRD);
      $finish;
    end

    if ((TXPCSRESET_TIME >= 5'b00000) && (TXPCSRESET_TIME <= 5'b11111))
      TXPCSRESET_TIME_BINARY = TXPCSRESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute TXPCSRESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TXPCSRESET_TIME);
      $finish;
    end

    if ((TXPH_MONITOR_SEL >= 5'b00000) && (TXPH_MONITOR_SEL <= 5'b11111))
      TXPH_MONITOR_SEL_BINARY = TXPH_MONITOR_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute TXPH_MONITOR_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TXPH_MONITOR_SEL);
      $finish;
    end

    if ((TXPMARESET_TIME >= 5'b00000) && (TXPMARESET_TIME <= 5'b11111))
      TXPMARESET_TIME_BINARY = TXPMARESET_TIME;
    else begin
      $display("Attribute Syntax Error : The Attribute TXPMARESET_TIME on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TXPMARESET_TIME);
      $finish;
    end

    if ((TX_CLKMUX_PD >= 1'b0) && (TX_CLKMUX_PD <= 1'b1))
      TX_CLKMUX_PD_BINARY = TX_CLKMUX_PD;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_CLKMUX_PD on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", TX_CLKMUX_PD);
      $finish;
    end

    if ((TX_DEEMPH0 >= 5'b00000) && (TX_DEEMPH0 <= 5'b11111))
      TX_DEEMPH0_BINARY = TX_DEEMPH0;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_DEEMPH0 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TX_DEEMPH0);
      $finish;
    end

    if ((TX_DEEMPH1 >= 5'b00000) && (TX_DEEMPH1 <= 5'b11111))
      TX_DEEMPH1_BINARY = TX_DEEMPH1;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_DEEMPH1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 5'b00000 to 5'b11111.", TX_DEEMPH1);
      $finish;
    end

    if ((TX_EIDLE_ASSERT_DELAY >= 3'b000) && (TX_EIDLE_ASSERT_DELAY <= 3'b111))
      TX_EIDLE_ASSERT_DELAY_BINARY = TX_EIDLE_ASSERT_DELAY;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_EIDLE_ASSERT_DELAY on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", TX_EIDLE_ASSERT_DELAY);
      $finish;
    end

    if ((TX_EIDLE_DEASSERT_DELAY >= 3'b000) && (TX_EIDLE_DEASSERT_DELAY <= 3'b111))
      TX_EIDLE_DEASSERT_DELAY_BINARY = TX_EIDLE_DEASSERT_DELAY;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_EIDLE_DEASSERT_DELAY on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", TX_EIDLE_DEASSERT_DELAY);
      $finish;
    end

    if ((TX_INT_DATAWIDTH >= 0) && (TX_INT_DATAWIDTH <= 1))
      TX_INT_DATAWIDTH_BINARY = TX_INT_DATAWIDTH;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_INT_DATAWIDTH on X_GTXE2_CHANNEL instance %m is set to %d.  Legal values for this attribute are  0 to 1.", TX_INT_DATAWIDTH);
      $finish;
    end

    if ((TX_MAINCURSOR_SEL >= 1'b0) && (TX_MAINCURSOR_SEL <= 1'b1))
      TX_MAINCURSOR_SEL_BINARY = TX_MAINCURSOR_SEL;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MAINCURSOR_SEL on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", TX_MAINCURSOR_SEL);
      $finish;
    end

    if ((TX_MARGIN_FULL_0 >= 7'b0000000) && (TX_MARGIN_FULL_0 <= 7'b1111111))
      TX_MARGIN_FULL_0_BINARY = TX_MARGIN_FULL_0;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_FULL_0 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_FULL_0);
      $finish;
    end

    if ((TX_MARGIN_FULL_1 >= 7'b0000000) && (TX_MARGIN_FULL_1 <= 7'b1111111))
      TX_MARGIN_FULL_1_BINARY = TX_MARGIN_FULL_1;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_FULL_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_FULL_1);
      $finish;
    end

    if ((TX_MARGIN_FULL_2 >= 7'b0000000) && (TX_MARGIN_FULL_2 <= 7'b1111111))
      TX_MARGIN_FULL_2_BINARY = TX_MARGIN_FULL_2;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_FULL_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_FULL_2);
      $finish;
    end

    if ((TX_MARGIN_FULL_3 >= 7'b0000000) && (TX_MARGIN_FULL_3 <= 7'b1111111))
      TX_MARGIN_FULL_3_BINARY = TX_MARGIN_FULL_3;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_FULL_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_FULL_3);
      $finish;
    end

    if ((TX_MARGIN_FULL_4 >= 7'b0000000) && (TX_MARGIN_FULL_4 <= 7'b1111111))
      TX_MARGIN_FULL_4_BINARY = TX_MARGIN_FULL_4;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_FULL_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_FULL_4);
      $finish;
    end

    if ((TX_MARGIN_LOW_0 >= 7'b0000000) && (TX_MARGIN_LOW_0 <= 7'b1111111))
      TX_MARGIN_LOW_0_BINARY = TX_MARGIN_LOW_0;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_LOW_0 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_LOW_0);
      $finish;
    end

    if ((TX_MARGIN_LOW_1 >= 7'b0000000) && (TX_MARGIN_LOW_1 <= 7'b1111111))
      TX_MARGIN_LOW_1_BINARY = TX_MARGIN_LOW_1;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_LOW_1 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_LOW_1);
      $finish;
    end

    if ((TX_MARGIN_LOW_2 >= 7'b0000000) && (TX_MARGIN_LOW_2 <= 7'b1111111))
      TX_MARGIN_LOW_2_BINARY = TX_MARGIN_LOW_2;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_LOW_2 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_LOW_2);
      $finish;
    end

    if ((TX_MARGIN_LOW_3 >= 7'b0000000) && (TX_MARGIN_LOW_3 <= 7'b1111111))
      TX_MARGIN_LOW_3_BINARY = TX_MARGIN_LOW_3;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_LOW_3 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_LOW_3);
      $finish;
    end

    if ((TX_MARGIN_LOW_4 >= 7'b0000000) && (TX_MARGIN_LOW_4 <= 7'b1111111))
      TX_MARGIN_LOW_4_BINARY = TX_MARGIN_LOW_4;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_MARGIN_LOW_4 on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 7'b0000000 to 7'b1111111.", TX_MARGIN_LOW_4);
      $finish;
    end

    if ((TX_PREDRIVER_MODE >= 1'b0) && (TX_PREDRIVER_MODE <= 1'b1))
      TX_PREDRIVER_MODE_BINARY = TX_PREDRIVER_MODE;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_PREDRIVER_MODE on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", TX_PREDRIVER_MODE);
      $finish;
    end

    if ((TX_QPI_STATUS_EN >= 1'b0) && (TX_QPI_STATUS_EN <= 1'b1))
      TX_QPI_STATUS_EN_BINARY = TX_QPI_STATUS_EN;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_QPI_STATUS_EN on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", TX_QPI_STATUS_EN);
      $finish;
    end

    if ((TX_RXDETECT_REF >= 3'b000) && (TX_RXDETECT_REF <= 3'b111))
      TX_RXDETECT_REF_BINARY = TX_RXDETECT_REF;
    else begin
      $display("Attribute Syntax Error : The Attribute TX_RXDETECT_REF on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 3'b000 to 3'b111.", TX_RXDETECT_REF);
      $finish;
    end

    if ((UCODEER_CLR >= 1'b0) && (UCODEER_CLR <= 1'b1))
      UCODEER_CLR_BINARY = UCODEER_CLR;
    else begin
      $display("Attribute Syntax Error : The Attribute UCODEER_CLR on X_GTXE2_CHANNEL instance %m is set to %b.  Legal values for this attribute are 1'b0 to 1'b1.", UCODEER_CLR);
      $finish;
    end

  end

  buf B_CPLLFBCLKLOST (CPLLFBCLKLOST, CPLLFBCLKLOST_OUT);
  buf B_CPLLLOCK (CPLLLOCK, CPLLLOCK_OUT);
  buf B_CPLLREFCLKLOST (CPLLREFCLKLOST, CPLLREFCLKLOST_OUT);
  buf B_DMONITOROUT0 (DMONITOROUT[0], DMONITOROUT_OUT[0]);
  buf B_DMONITOROUT1 (DMONITOROUT[1], DMONITOROUT_OUT[1]);
  buf B_DMONITOROUT2 (DMONITOROUT[2], DMONITOROUT_OUT[2]);
  buf B_DMONITOROUT3 (DMONITOROUT[3], DMONITOROUT_OUT[3]);
  buf B_DMONITOROUT4 (DMONITOROUT[4], DMONITOROUT_OUT[4]);
  buf B_DMONITOROUT5 (DMONITOROUT[5], DMONITOROUT_OUT[5]);
  buf B_DMONITOROUT6 (DMONITOROUT[6], DMONITOROUT_OUT[6]);
  buf B_DMONITOROUT7 (DMONITOROUT[7], DMONITOROUT_OUT[7]);
  buf B_DRPDO0 (DRPDO[0], DRPDO_OUT[0]);
  buf B_DRPDO1 (DRPDO[1], DRPDO_OUT[1]);
  buf B_DRPDO10 (DRPDO[10], DRPDO_OUT[10]);
  buf B_DRPDO11 (DRPDO[11], DRPDO_OUT[11]);
  buf B_DRPDO12 (DRPDO[12], DRPDO_OUT[12]);
  buf B_DRPDO13 (DRPDO[13], DRPDO_OUT[13]);
  buf B_DRPDO14 (DRPDO[14], DRPDO_OUT[14]);
  buf B_DRPDO15 (DRPDO[15], DRPDO_OUT[15]);
  buf B_DRPDO2 (DRPDO[2], DRPDO_OUT[2]);
  buf B_DRPDO3 (DRPDO[3], DRPDO_OUT[3]);
  buf B_DRPDO4 (DRPDO[4], DRPDO_OUT[4]);
  buf B_DRPDO5 (DRPDO[5], DRPDO_OUT[5]);
  buf B_DRPDO6 (DRPDO[6], DRPDO_OUT[6]);
  buf B_DRPDO7 (DRPDO[7], DRPDO_OUT[7]);
  buf B_DRPDO8 (DRPDO[8], DRPDO_OUT[8]);
  buf B_DRPDO9 (DRPDO[9], DRPDO_OUT[9]);
  buf B_DRPRDY (DRPRDY, DRPRDY_OUT);
  buf B_EYESCANDATAERROR (EYESCANDATAERROR, EYESCANDATAERROR_OUT);
  buf B_GTREFCLKMONITOR (GTREFCLKMONITOR, GTREFCLKMONITOR_OUT);
  buf B_GTXTXN (GTXTXN, GTXTXN_OUT);
  buf B_GTXTXP (GTXTXP, GTXTXP_OUT);
  buf B_PCSRSVDOUT0 (PCSRSVDOUT[0], PCSRSVDOUT_OUT[0]);
  buf B_PCSRSVDOUT1 (PCSRSVDOUT[1], PCSRSVDOUT_OUT[1]);
  buf B_PCSRSVDOUT10 (PCSRSVDOUT[10], PCSRSVDOUT_OUT[10]);
  buf B_PCSRSVDOUT11 (PCSRSVDOUT[11], PCSRSVDOUT_OUT[11]);
  buf B_PCSRSVDOUT12 (PCSRSVDOUT[12], PCSRSVDOUT_OUT[12]);
  buf B_PCSRSVDOUT13 (PCSRSVDOUT[13], PCSRSVDOUT_OUT[13]);
  buf B_PCSRSVDOUT14 (PCSRSVDOUT[14], PCSRSVDOUT_OUT[14]);
  buf B_PCSRSVDOUT15 (PCSRSVDOUT[15], PCSRSVDOUT_OUT[15]);
  buf B_PCSRSVDOUT2 (PCSRSVDOUT[2], PCSRSVDOUT_OUT[2]);
  buf B_PCSRSVDOUT3 (PCSRSVDOUT[3], PCSRSVDOUT_OUT[3]);
  buf B_PCSRSVDOUT4 (PCSRSVDOUT[4], PCSRSVDOUT_OUT[4]);
  buf B_PCSRSVDOUT5 (PCSRSVDOUT[5], PCSRSVDOUT_OUT[5]);
  buf B_PCSRSVDOUT6 (PCSRSVDOUT[6], PCSRSVDOUT_OUT[6]);
  buf B_PCSRSVDOUT7 (PCSRSVDOUT[7], PCSRSVDOUT_OUT[7]);
  buf B_PCSRSVDOUT8 (PCSRSVDOUT[8], PCSRSVDOUT_OUT[8]);
  buf B_PCSRSVDOUT9 (PCSRSVDOUT[9], PCSRSVDOUT_OUT[9]);
  buf B_PHYSTATUS (PHYSTATUS, PHYSTATUS_OUT);
  buf B_RXBUFSTATUS0 (RXBUFSTATUS[0], RXBUFSTATUS_OUT[0]);
  buf B_RXBUFSTATUS1 (RXBUFSTATUS[1], RXBUFSTATUS_OUT[1]);
  buf B_RXBUFSTATUS2 (RXBUFSTATUS[2], RXBUFSTATUS_OUT[2]);
  buf B_RXBYTEISALIGNED (RXBYTEISALIGNED, RXBYTEISALIGNED_OUT);
  buf B_RXBYTEREALIGN (RXBYTEREALIGN, RXBYTEREALIGN_OUT);
  buf B_RXCDRLOCK (RXCDRLOCK, RXCDRLOCK_OUT);
  buf B_RXCHANBONDSEQ (RXCHANBONDSEQ, RXCHANBONDSEQ_OUT);
  buf B_RXCHANISALIGNED (RXCHANISALIGNED, RXCHANISALIGNED_OUT);
  buf B_RXCHANREALIGN (RXCHANREALIGN, RXCHANREALIGN_OUT);
  buf B_RXCHARISCOMMA0 (RXCHARISCOMMA[0], RXCHARISCOMMA_OUT[0]);
  buf B_RXCHARISCOMMA1 (RXCHARISCOMMA[1], RXCHARISCOMMA_OUT[1]);
  buf B_RXCHARISCOMMA2 (RXCHARISCOMMA[2], RXCHARISCOMMA_OUT[2]);
  buf B_RXCHARISCOMMA3 (RXCHARISCOMMA[3], RXCHARISCOMMA_OUT[3]);
  buf B_RXCHARISCOMMA4 (RXCHARISCOMMA[4], RXCHARISCOMMA_OUT[4]);
  buf B_RXCHARISCOMMA5 (RXCHARISCOMMA[5], RXCHARISCOMMA_OUT[5]);
  buf B_RXCHARISCOMMA6 (RXCHARISCOMMA[6], RXCHARISCOMMA_OUT[6]);
  buf B_RXCHARISCOMMA7 (RXCHARISCOMMA[7], RXCHARISCOMMA_OUT[7]);
  buf B_RXCHARISK0 (RXCHARISK[0], RXCHARISK_OUT[0]);
  buf B_RXCHARISK1 (RXCHARISK[1], RXCHARISK_OUT[1]);
  buf B_RXCHARISK2 (RXCHARISK[2], RXCHARISK_OUT[2]);
  buf B_RXCHARISK3 (RXCHARISK[3], RXCHARISK_OUT[3]);
  buf B_RXCHARISK4 (RXCHARISK[4], RXCHARISK_OUT[4]);
  buf B_RXCHARISK5 (RXCHARISK[5], RXCHARISK_OUT[5]);
  buf B_RXCHARISK6 (RXCHARISK[6], RXCHARISK_OUT[6]);
  buf B_RXCHARISK7 (RXCHARISK[7], RXCHARISK_OUT[7]);
  buf B_RXCHBONDO0 (RXCHBONDO[0], RXCHBONDO_OUT[0]);
  buf B_RXCHBONDO1 (RXCHBONDO[1], RXCHBONDO_OUT[1]);
  buf B_RXCHBONDO2 (RXCHBONDO[2], RXCHBONDO_OUT[2]);
  buf B_RXCHBONDO3 (RXCHBONDO[3], RXCHBONDO_OUT[3]);
  buf B_RXCHBONDO4 (RXCHBONDO[4], RXCHBONDO_OUT[4]);
  buf B_RXCLKCORCNT0 (RXCLKCORCNT[0], RXCLKCORCNT_OUT[0]);
  buf B_RXCLKCORCNT1 (RXCLKCORCNT[1], RXCLKCORCNT_OUT[1]);
  buf B_RXCOMINITDET (RXCOMINITDET, RXCOMINITDET_OUT);
  buf B_RXCOMMADET (RXCOMMADET, RXCOMMADET_OUT);
  buf B_RXCOMSASDET (RXCOMSASDET, RXCOMSASDET_OUT);
  buf B_RXCOMWAKEDET (RXCOMWAKEDET, RXCOMWAKEDET_OUT);
  buf B_RXDATA0 (RXDATA[0], RXDATA_OUT[0]);
  buf B_RXDATA1 (RXDATA[1], RXDATA_OUT[1]);
  buf B_RXDATA10 (RXDATA[10], RXDATA_OUT[10]);
  buf B_RXDATA11 (RXDATA[11], RXDATA_OUT[11]);
  buf B_RXDATA12 (RXDATA[12], RXDATA_OUT[12]);
  buf B_RXDATA13 (RXDATA[13], RXDATA_OUT[13]);
  buf B_RXDATA14 (RXDATA[14], RXDATA_OUT[14]);
  buf B_RXDATA15 (RXDATA[15], RXDATA_OUT[15]);
  buf B_RXDATA16 (RXDATA[16], RXDATA_OUT[16]);
  buf B_RXDATA17 (RXDATA[17], RXDATA_OUT[17]);
  buf B_RXDATA18 (RXDATA[18], RXDATA_OUT[18]);
  buf B_RXDATA19 (RXDATA[19], RXDATA_OUT[19]);
  buf B_RXDATA2 (RXDATA[2], RXDATA_OUT[2]);
  buf B_RXDATA20 (RXDATA[20], RXDATA_OUT[20]);
  buf B_RXDATA21 (RXDATA[21], RXDATA_OUT[21]);
  buf B_RXDATA22 (RXDATA[22], RXDATA_OUT[22]);
  buf B_RXDATA23 (RXDATA[23], RXDATA_OUT[23]);
  buf B_RXDATA24 (RXDATA[24], RXDATA_OUT[24]);
  buf B_RXDATA25 (RXDATA[25], RXDATA_OUT[25]);
  buf B_RXDATA26 (RXDATA[26], RXDATA_OUT[26]);
  buf B_RXDATA27 (RXDATA[27], RXDATA_OUT[27]);
  buf B_RXDATA28 (RXDATA[28], RXDATA_OUT[28]);
  buf B_RXDATA29 (RXDATA[29], RXDATA_OUT[29]);
  buf B_RXDATA3 (RXDATA[3], RXDATA_OUT[3]);
  buf B_RXDATA30 (RXDATA[30], RXDATA_OUT[30]);
  buf B_RXDATA31 (RXDATA[31], RXDATA_OUT[31]);
  buf B_RXDATA32 (RXDATA[32], RXDATA_OUT[32]);
  buf B_RXDATA33 (RXDATA[33], RXDATA_OUT[33]);
  buf B_RXDATA34 (RXDATA[34], RXDATA_OUT[34]);
  buf B_RXDATA35 (RXDATA[35], RXDATA_OUT[35]);
  buf B_RXDATA36 (RXDATA[36], RXDATA_OUT[36]);
  buf B_RXDATA37 (RXDATA[37], RXDATA_OUT[37]);
  buf B_RXDATA38 (RXDATA[38], RXDATA_OUT[38]);
  buf B_RXDATA39 (RXDATA[39], RXDATA_OUT[39]);
  buf B_RXDATA4 (RXDATA[4], RXDATA_OUT[4]);
  buf B_RXDATA40 (RXDATA[40], RXDATA_OUT[40]);
  buf B_RXDATA41 (RXDATA[41], RXDATA_OUT[41]);
  buf B_RXDATA42 (RXDATA[42], RXDATA_OUT[42]);
  buf B_RXDATA43 (RXDATA[43], RXDATA_OUT[43]);
  buf B_RXDATA44 (RXDATA[44], RXDATA_OUT[44]);
  buf B_RXDATA45 (RXDATA[45], RXDATA_OUT[45]);
  buf B_RXDATA46 (RXDATA[46], RXDATA_OUT[46]);
  buf B_RXDATA47 (RXDATA[47], RXDATA_OUT[47]);
  buf B_RXDATA48 (RXDATA[48], RXDATA_OUT[48]);
  buf B_RXDATA49 (RXDATA[49], RXDATA_OUT[49]);
  buf B_RXDATA5 (RXDATA[5], RXDATA_OUT[5]);
  buf B_RXDATA50 (RXDATA[50], RXDATA_OUT[50]);
  buf B_RXDATA51 (RXDATA[51], RXDATA_OUT[51]);
  buf B_RXDATA52 (RXDATA[52], RXDATA_OUT[52]);
  buf B_RXDATA53 (RXDATA[53], RXDATA_OUT[53]);
  buf B_RXDATA54 (RXDATA[54], RXDATA_OUT[54]);
  buf B_RXDATA55 (RXDATA[55], RXDATA_OUT[55]);
  buf B_RXDATA56 (RXDATA[56], RXDATA_OUT[56]);
  buf B_RXDATA57 (RXDATA[57], RXDATA_OUT[57]);
  buf B_RXDATA58 (RXDATA[58], RXDATA_OUT[58]);
  buf B_RXDATA59 (RXDATA[59], RXDATA_OUT[59]);
  buf B_RXDATA6 (RXDATA[6], RXDATA_OUT[6]);
  buf B_RXDATA60 (RXDATA[60], RXDATA_OUT[60]);
  buf B_RXDATA61 (RXDATA[61], RXDATA_OUT[61]);
  buf B_RXDATA62 (RXDATA[62], RXDATA_OUT[62]);
  buf B_RXDATA63 (RXDATA[63], RXDATA_OUT[63]);
  buf B_RXDATA7 (RXDATA[7], RXDATA_OUT[7]);
  buf B_RXDATA8 (RXDATA[8], RXDATA_OUT[8]);
  buf B_RXDATA9 (RXDATA[9], RXDATA_OUT[9]);
  buf B_RXDATAVALID (RXDATAVALID, RXDATAVALID_OUT);
  buf B_RXDISPERR0 (RXDISPERR[0], RXDISPERR_OUT[0]);
  buf B_RXDISPERR1 (RXDISPERR[1], RXDISPERR_OUT[1]);
  buf B_RXDISPERR2 (RXDISPERR[2], RXDISPERR_OUT[2]);
  buf B_RXDISPERR3 (RXDISPERR[3], RXDISPERR_OUT[3]);
  buf B_RXDISPERR4 (RXDISPERR[4], RXDISPERR_OUT[4]);
  buf B_RXDISPERR5 (RXDISPERR[5], RXDISPERR_OUT[5]);
  buf B_RXDISPERR6 (RXDISPERR[6], RXDISPERR_OUT[6]);
  buf B_RXDISPERR7 (RXDISPERR[7], RXDISPERR_OUT[7]);
  buf B_RXDLYSRESETDONE (RXDLYSRESETDONE, RXDLYSRESETDONE_OUT);
  buf B_RXELECIDLE (RXELECIDLE, RXELECIDLE_OUT);
  buf B_RXHEADER0 (RXHEADER[0], RXHEADER_OUT[0]);
  buf B_RXHEADER1 (RXHEADER[1], RXHEADER_OUT[1]);
  buf B_RXHEADER2 (RXHEADER[2], RXHEADER_OUT[2]);
  buf B_RXHEADERVALID (RXHEADERVALID, RXHEADERVALID_OUT);
  buf B_RXMONITOROUT0 (RXMONITOROUT[0], RXMONITOROUT_OUT[0]);
  buf B_RXMONITOROUT1 (RXMONITOROUT[1], RXMONITOROUT_OUT[1]);
  buf B_RXMONITOROUT2 (RXMONITOROUT[2], RXMONITOROUT_OUT[2]);
  buf B_RXMONITOROUT3 (RXMONITOROUT[3], RXMONITOROUT_OUT[3]);
  buf B_RXMONITOROUT4 (RXMONITOROUT[4], RXMONITOROUT_OUT[4]);
  buf B_RXMONITOROUT5 (RXMONITOROUT[5], RXMONITOROUT_OUT[5]);
  buf B_RXMONITOROUT6 (RXMONITOROUT[6], RXMONITOROUT_OUT[6]);
  buf B_RXNOTINTABLE0 (RXNOTINTABLE[0], RXNOTINTABLE_OUT[0]);
  buf B_RXNOTINTABLE1 (RXNOTINTABLE[1], RXNOTINTABLE_OUT[1]);
  buf B_RXNOTINTABLE2 (RXNOTINTABLE[2], RXNOTINTABLE_OUT[2]);
  buf B_RXNOTINTABLE3 (RXNOTINTABLE[3], RXNOTINTABLE_OUT[3]);
  buf B_RXNOTINTABLE4 (RXNOTINTABLE[4], RXNOTINTABLE_OUT[4]);
  buf B_RXNOTINTABLE5 (RXNOTINTABLE[5], RXNOTINTABLE_OUT[5]);
  buf B_RXNOTINTABLE6 (RXNOTINTABLE[6], RXNOTINTABLE_OUT[6]);
  buf B_RXNOTINTABLE7 (RXNOTINTABLE[7], RXNOTINTABLE_OUT[7]);
  buf B_RXOUTCLK (RXOUTCLK, RXOUTCLK_OUT);
  buf B_RXOUTCLKFABRIC (RXOUTCLKFABRIC, RXOUTCLKFABRIC_OUT);
  buf B_RXOUTCLKPCS (RXOUTCLKPCS, RXOUTCLKPCS_OUT);
  buf B_RXPHALIGNDONE (RXPHALIGNDONE, RXPHALIGNDONE_OUT);
  buf B_RXPHMONITOR0 (RXPHMONITOR[0], RXPHMONITOR_OUT[0]);
  buf B_RXPHMONITOR1 (RXPHMONITOR[1], RXPHMONITOR_OUT[1]);
  buf B_RXPHMONITOR2 (RXPHMONITOR[2], RXPHMONITOR_OUT[2]);
  buf B_RXPHMONITOR3 (RXPHMONITOR[3], RXPHMONITOR_OUT[3]);
  buf B_RXPHMONITOR4 (RXPHMONITOR[4], RXPHMONITOR_OUT[4]);
  buf B_RXPHSLIPMONITOR0 (RXPHSLIPMONITOR[0], RXPHSLIPMONITOR_OUT[0]);
  buf B_RXPHSLIPMONITOR1 (RXPHSLIPMONITOR[1], RXPHSLIPMONITOR_OUT[1]);
  buf B_RXPHSLIPMONITOR2 (RXPHSLIPMONITOR[2], RXPHSLIPMONITOR_OUT[2]);
  buf B_RXPHSLIPMONITOR3 (RXPHSLIPMONITOR[3], RXPHSLIPMONITOR_OUT[3]);
  buf B_RXPHSLIPMONITOR4 (RXPHSLIPMONITOR[4], RXPHSLIPMONITOR_OUT[4]);
  buf B_RXPRBSERR (RXPRBSERR, RXPRBSERR_OUT);
  buf B_RXQPISENN (RXQPISENN, RXQPISENN_OUT);
  buf B_RXQPISENP (RXQPISENP, RXQPISENP_OUT);
  buf B_RXRATEDONE (RXRATEDONE, RXRATEDONE_OUT);
  buf B_RXRESETDONE (RXRESETDONE, RXRESETDONE_OUT);
  buf B_RXSTARTOFSEQ (RXSTARTOFSEQ, RXSTARTOFSEQ_OUT);
  buf B_RXSTATUS0 (RXSTATUS[0], RXSTATUS_OUT[0]);
  buf B_RXSTATUS1 (RXSTATUS[1], RXSTATUS_OUT[1]);
  buf B_RXSTATUS2 (RXSTATUS[2], RXSTATUS_OUT[2]);
  buf B_RXVALID (RXVALID, RXVALID_OUT);
  buf B_TSTOUT0 (TSTOUT[0], TSTOUT_OUT[0]);
  buf B_TSTOUT1 (TSTOUT[1], TSTOUT_OUT[1]);
  buf B_TSTOUT2 (TSTOUT[2], TSTOUT_OUT[2]);
  buf B_TSTOUT3 (TSTOUT[3], TSTOUT_OUT[3]);
  buf B_TSTOUT4 (TSTOUT[4], TSTOUT_OUT[4]);
  buf B_TSTOUT5 (TSTOUT[5], TSTOUT_OUT[5]);
  buf B_TSTOUT6 (TSTOUT[6], TSTOUT_OUT[6]);
  buf B_TSTOUT7 (TSTOUT[7], TSTOUT_OUT[7]);
  buf B_TSTOUT8 (TSTOUT[8], TSTOUT_OUT[8]);
  buf B_TSTOUT9 (TSTOUT[9], TSTOUT_OUT[9]);
  buf B_TXBUFSTATUS0 (TXBUFSTATUS[0], TXBUFSTATUS_OUT[0]);
  buf B_TXBUFSTATUS1 (TXBUFSTATUS[1], TXBUFSTATUS_OUT[1]);
  buf B_TXCOMFINISH (TXCOMFINISH, TXCOMFINISH_OUT);
  buf B_TXDLYSRESETDONE (TXDLYSRESETDONE, TXDLYSRESETDONE_OUT);
  buf B_TXGEARBOXREADY (TXGEARBOXREADY, TXGEARBOXREADY_OUT);
  buf B_TXOUTCLK (TXOUTCLK, TXOUTCLK_OUT);
  buf B_TXOUTCLKFABRIC (TXOUTCLKFABRIC, TXOUTCLKFABRIC_OUT);
  buf B_TXOUTCLKPCS (TXOUTCLKPCS, TXOUTCLKPCS_OUT);
  buf B_TXPHALIGNDONE (TXPHALIGNDONE, TXPHALIGNDONE_OUT);
  buf B_TXPHINITDONE (TXPHINITDONE, TXPHINITDONE_OUT);
  buf B_TXQPISENN (TXQPISENN, TXQPISENN_OUT);
  buf B_TXQPISENP (TXQPISENP, TXQPISENP_OUT);
  buf B_TXRATEDONE (TXRATEDONE, TXRATEDONE_OUT);
  buf B_TXRESETDONE (TXRESETDONE, TXRESETDONE_OUT);

  buf B_CFGRESET (CFGRESET_IN, CFGRESET);
  buf B_CLKRSVD0 (CLKRSVD_IN[0], CLKRSVD[0]);
  buf B_CLKRSVD1 (CLKRSVD_IN[1], CLKRSVD[1]);
  buf B_CLKRSVD2 (CLKRSVD_IN[2], CLKRSVD[2]);
  buf B_CLKRSVD3 (CLKRSVD_IN[3], CLKRSVD[3]);
  buf B_CPLLLOCKDETCLK (CPLLLOCKDETCLK_IN, CPLLLOCKDETCLK);
  buf B_CPLLLOCKEN (CPLLLOCKEN_IN, CPLLLOCKEN);
  buf B_CPLLPD (CPLLPD_IN, CPLLPD);
  buf B_CPLLREFCLKSEL0 (CPLLREFCLKSEL_IN[0], CPLLREFCLKSEL[0]);
  buf B_CPLLREFCLKSEL1 (CPLLREFCLKSEL_IN[1], CPLLREFCLKSEL[1]);
  buf B_CPLLREFCLKSEL2 (CPLLREFCLKSEL_IN[2], CPLLREFCLKSEL[2]);
  buf B_CPLLRESET (CPLLRESET_IN, CPLLRESET);
  buf B_DRPADDR0 (DRPADDR_IN[0], DRPADDR[0]);
  buf B_DRPADDR1 (DRPADDR_IN[1], DRPADDR[1]);
  buf B_DRPADDR2 (DRPADDR_IN[2], DRPADDR[2]);
  buf B_DRPADDR3 (DRPADDR_IN[3], DRPADDR[3]);
  buf B_DRPADDR4 (DRPADDR_IN[4], DRPADDR[4]);
  buf B_DRPADDR5 (DRPADDR_IN[5], DRPADDR[5]);
  buf B_DRPADDR6 (DRPADDR_IN[6], DRPADDR[6]);
  buf B_DRPADDR7 (DRPADDR_IN[7], DRPADDR[7]);
  buf B_DRPADDR8 (DRPADDR_IN[8], DRPADDR[8]);
  buf B_DRPCLK (DRPCLK_IN, DRPCLK);
  buf B_DRPDI0 (DRPDI_IN[0], DRPDI[0]);
  buf B_DRPDI1 (DRPDI_IN[1], DRPDI[1]);
  buf B_DRPDI10 (DRPDI_IN[10], DRPDI[10]);
  buf B_DRPDI11 (DRPDI_IN[11], DRPDI[11]);
  buf B_DRPDI12 (DRPDI_IN[12], DRPDI[12]);
  buf B_DRPDI13 (DRPDI_IN[13], DRPDI[13]);
  buf B_DRPDI14 (DRPDI_IN[14], DRPDI[14]);
  buf B_DRPDI15 (DRPDI_IN[15], DRPDI[15]);
  buf B_DRPDI2 (DRPDI_IN[2], DRPDI[2]);
  buf B_DRPDI3 (DRPDI_IN[3], DRPDI[3]);
  buf B_DRPDI4 (DRPDI_IN[4], DRPDI[4]);
  buf B_DRPDI5 (DRPDI_IN[5], DRPDI[5]);
  buf B_DRPDI6 (DRPDI_IN[6], DRPDI[6]);
  buf B_DRPDI7 (DRPDI_IN[7], DRPDI[7]);
  buf B_DRPDI8 (DRPDI_IN[8], DRPDI[8]);
  buf B_DRPDI9 (DRPDI_IN[9], DRPDI[9]);
  buf B_DRPEN (DRPEN_IN, DRPEN);
  buf B_DRPWE (DRPWE_IN, DRPWE);
  buf B_EYESCANMODE (EYESCANMODE_IN, EYESCANMODE);
  buf B_EYESCANRESET (EYESCANRESET_IN, EYESCANRESET);
  buf B_EYESCANTRIGGER (EYESCANTRIGGER_IN, EYESCANTRIGGER);
  buf B_GTGREFCLK (GTGREFCLK_IN, GTGREFCLK);
  buf B_GTNORTHREFCLK0 (GTNORTHREFCLK0_IN, GTNORTHREFCLK0);
  buf B_GTNORTHREFCLK1 (GTNORTHREFCLK1_IN, GTNORTHREFCLK1);
  buf B_GTREFCLK0 (GTREFCLK0_IN, GTREFCLK0);
  buf B_GTREFCLK1 (GTREFCLK1_IN, GTREFCLK1);
  buf B_GTRESETSEL (GTRESETSEL_IN, GTRESETSEL);
  buf B_GTRSVD0 (GTRSVD_IN[0], GTRSVD[0]);
  buf B_GTRSVD1 (GTRSVD_IN[1], GTRSVD[1]);
  buf B_GTRSVD10 (GTRSVD_IN[10], GTRSVD[10]);
  buf B_GTRSVD11 (GTRSVD_IN[11], GTRSVD[11]);
  buf B_GTRSVD12 (GTRSVD_IN[12], GTRSVD[12]);
  buf B_GTRSVD13 (GTRSVD_IN[13], GTRSVD[13]);
  buf B_GTRSVD14 (GTRSVD_IN[14], GTRSVD[14]);
  buf B_GTRSVD15 (GTRSVD_IN[15], GTRSVD[15]);
  buf B_GTRSVD2 (GTRSVD_IN[2], GTRSVD[2]);
  buf B_GTRSVD3 (GTRSVD_IN[3], GTRSVD[3]);
  buf B_GTRSVD4 (GTRSVD_IN[4], GTRSVD[4]);
  buf B_GTRSVD5 (GTRSVD_IN[5], GTRSVD[5]);
  buf B_GTRSVD6 (GTRSVD_IN[6], GTRSVD[6]);
  buf B_GTRSVD7 (GTRSVD_IN[7], GTRSVD[7]);
  buf B_GTRSVD8 (GTRSVD_IN[8], GTRSVD[8]);
  buf B_GTRSVD9 (GTRSVD_IN[9], GTRSVD[9]);
  buf B_GTRXRESET (GTRXRESET_IN, GTRXRESET);
  buf B_GTSOUTHREFCLK0 (GTSOUTHREFCLK0_IN, GTSOUTHREFCLK0);
  buf B_GTSOUTHREFCLK1 (GTSOUTHREFCLK1_IN, GTSOUTHREFCLK1);
  buf B_GTTXRESET (GTTXRESET_IN, GTTXRESET);
  buf B_GTXRXN (GTXRXN_IN, GTXRXN);
  buf B_GTXRXP (GTXRXP_IN, GTXRXP);
  buf B_LOOPBACK0 (LOOPBACK_IN[0], LOOPBACK[0]);
  buf B_LOOPBACK1 (LOOPBACK_IN[1], LOOPBACK[1]);
  buf B_LOOPBACK2 (LOOPBACK_IN[2], LOOPBACK[2]);
  buf B_PCSRSVDIN0 (PCSRSVDIN_IN[0], PCSRSVDIN[0]);
  buf B_PCSRSVDIN1 (PCSRSVDIN_IN[1], PCSRSVDIN[1]);
  buf B_PCSRSVDIN10 (PCSRSVDIN_IN[10], PCSRSVDIN[10]);
  buf B_PCSRSVDIN11 (PCSRSVDIN_IN[11], PCSRSVDIN[11]);
  buf B_PCSRSVDIN12 (PCSRSVDIN_IN[12], PCSRSVDIN[12]);
  buf B_PCSRSVDIN13 (PCSRSVDIN_IN[13], PCSRSVDIN[13]);
  buf B_PCSRSVDIN14 (PCSRSVDIN_IN[14], PCSRSVDIN[14]);
  buf B_PCSRSVDIN15 (PCSRSVDIN_IN[15], PCSRSVDIN[15]);
  buf B_PCSRSVDIN2 (PCSRSVDIN_IN[2], PCSRSVDIN[2]);
  buf B_PCSRSVDIN20 (PCSRSVDIN2_IN[0], PCSRSVDIN2[0]);
  buf B_PCSRSVDIN21 (PCSRSVDIN2_IN[1], PCSRSVDIN2[1]);
  buf B_PCSRSVDIN22 (PCSRSVDIN2_IN[2], PCSRSVDIN2[2]);
  buf B_PCSRSVDIN23 (PCSRSVDIN2_IN[3], PCSRSVDIN2[3]);
  buf B_PCSRSVDIN24 (PCSRSVDIN2_IN[4], PCSRSVDIN2[4]);
  buf B_PCSRSVDIN3 (PCSRSVDIN_IN[3], PCSRSVDIN[3]);
  buf B_PCSRSVDIN4 (PCSRSVDIN_IN[4], PCSRSVDIN[4]);
  buf B_PCSRSVDIN5 (PCSRSVDIN_IN[5], PCSRSVDIN[5]);
  buf B_PCSRSVDIN6 (PCSRSVDIN_IN[6], PCSRSVDIN[6]);
  buf B_PCSRSVDIN7 (PCSRSVDIN_IN[7], PCSRSVDIN[7]);
  buf B_PCSRSVDIN8 (PCSRSVDIN_IN[8], PCSRSVDIN[8]);
  buf B_PCSRSVDIN9 (PCSRSVDIN_IN[9], PCSRSVDIN[9]);
  buf B_PMARSVDIN0 (PMARSVDIN_IN[0], PMARSVDIN[0]);
  buf B_PMARSVDIN1 (PMARSVDIN_IN[1], PMARSVDIN[1]);
  buf B_PMARSVDIN2 (PMARSVDIN_IN[2], PMARSVDIN[2]);
  buf B_PMARSVDIN20 (PMARSVDIN2_IN[0], PMARSVDIN2[0]);
  buf B_PMARSVDIN21 (PMARSVDIN2_IN[1], PMARSVDIN2[1]);
  buf B_PMARSVDIN22 (PMARSVDIN2_IN[2], PMARSVDIN2[2]);
  buf B_PMARSVDIN23 (PMARSVDIN2_IN[3], PMARSVDIN2[3]);
  buf B_PMARSVDIN24 (PMARSVDIN2_IN[4], PMARSVDIN2[4]);
  buf B_PMARSVDIN3 (PMARSVDIN_IN[3], PMARSVDIN[3]);
  buf B_PMARSVDIN4 (PMARSVDIN_IN[4], PMARSVDIN[4]);
  buf B_QPLLCLK (QPLLCLK_IN, QPLLCLK);
  buf B_QPLLREFCLK (QPLLREFCLK_IN, QPLLREFCLK);
  buf B_RESETOVRD (RESETOVRD_IN, RESETOVRD);
  buf B_RX8B10BEN (RX8B10BEN_IN, RX8B10BEN);
  buf B_RXBUFRESET (RXBUFRESET_IN, RXBUFRESET);
  buf B_RXCDRFREQRESET (RXCDRFREQRESET_IN, RXCDRFREQRESET);
  buf B_RXCDRHOLD (RXCDRHOLD_IN, RXCDRHOLD);
  buf B_RXCDROVRDEN (RXCDROVRDEN_IN, RXCDROVRDEN);
  buf B_RXCDRRESET (RXCDRRESET_IN, RXCDRRESET);
  buf B_RXCDRRESETRSV (RXCDRRESETRSV_IN, RXCDRRESETRSV);
  buf B_RXCHBONDEN (RXCHBONDEN_IN, RXCHBONDEN);
  buf B_RXCHBONDI0 (RXCHBONDI_IN[0], RXCHBONDI[0]);
  buf B_RXCHBONDI1 (RXCHBONDI_IN[1], RXCHBONDI[1]);
  buf B_RXCHBONDI2 (RXCHBONDI_IN[2], RXCHBONDI[2]);
  buf B_RXCHBONDI3 (RXCHBONDI_IN[3], RXCHBONDI[3]);
  buf B_RXCHBONDI4 (RXCHBONDI_IN[4], RXCHBONDI[4]);
  buf B_RXCHBONDLEVEL0 (RXCHBONDLEVEL_IN[0], RXCHBONDLEVEL[0]);
  buf B_RXCHBONDLEVEL1 (RXCHBONDLEVEL_IN[1], RXCHBONDLEVEL[1]);
  buf B_RXCHBONDLEVEL2 (RXCHBONDLEVEL_IN[2], RXCHBONDLEVEL[2]);
  buf B_RXCHBONDMASTER (RXCHBONDMASTER_IN, RXCHBONDMASTER);
  buf B_RXCHBONDSLAVE (RXCHBONDSLAVE_IN, RXCHBONDSLAVE);
  buf B_RXCOMMADETEN (RXCOMMADETEN_IN, RXCOMMADETEN);
  buf B_RXDDIEN (RXDDIEN_IN, RXDDIEN);
  buf B_RXDFEAGCHOLD (RXDFEAGCHOLD_IN, RXDFEAGCHOLD);
  buf B_RXDFEAGCOVRDEN (RXDFEAGCOVRDEN_IN, RXDFEAGCOVRDEN);
  buf B_RXDFECM1EN (RXDFECM1EN_IN, RXDFECM1EN);
  buf B_RXDFELFHOLD (RXDFELFHOLD_IN, RXDFELFHOLD);
  buf B_RXDFELFOVRDEN (RXDFELFOVRDEN_IN, RXDFELFOVRDEN);
  buf B_RXDFELPMRESET (RXDFELPMRESET_IN, RXDFELPMRESET);
  buf B_RXDFETAP2HOLD (RXDFETAP2HOLD_IN, RXDFETAP2HOLD);
  buf B_RXDFETAP2OVRDEN (RXDFETAP2OVRDEN_IN, RXDFETAP2OVRDEN);
  buf B_RXDFETAP3HOLD (RXDFETAP3HOLD_IN, RXDFETAP3HOLD);
  buf B_RXDFETAP3OVRDEN (RXDFETAP3OVRDEN_IN, RXDFETAP3OVRDEN);
  buf B_RXDFETAP4HOLD (RXDFETAP4HOLD_IN, RXDFETAP4HOLD);
  buf B_RXDFETAP4OVRDEN (RXDFETAP4OVRDEN_IN, RXDFETAP4OVRDEN);
  buf B_RXDFETAP5HOLD (RXDFETAP5HOLD_IN, RXDFETAP5HOLD);
  buf B_RXDFETAP5OVRDEN (RXDFETAP5OVRDEN_IN, RXDFETAP5OVRDEN);
  buf B_RXDFEUTHOLD (RXDFEUTHOLD_IN, RXDFEUTHOLD);
  buf B_RXDFEUTOVRDEN (RXDFEUTOVRDEN_IN, RXDFEUTOVRDEN);
  buf B_RXDFEVPHOLD (RXDFEVPHOLD_IN, RXDFEVPHOLD);
  buf B_RXDFEVPOVRDEN (RXDFEVPOVRDEN_IN, RXDFEVPOVRDEN);
  buf B_RXDFEVSEN (RXDFEVSEN_IN, RXDFEVSEN);
  buf B_RXDFEXYDEN (RXDFEXYDEN_IN, RXDFEXYDEN);
  buf B_RXDFEXYDHOLD (RXDFEXYDHOLD_IN, RXDFEXYDHOLD);
  buf B_RXDFEXYDOVRDEN (RXDFEXYDOVRDEN_IN, RXDFEXYDOVRDEN);
  buf B_RXDLYBYPASS (RXDLYBYPASS_IN, RXDLYBYPASS);
  buf B_RXDLYEN (RXDLYEN_IN, RXDLYEN);
  buf B_RXDLYOVRDEN (RXDLYOVRDEN_IN, RXDLYOVRDEN);
  buf B_RXDLYSRESET (RXDLYSRESET_IN, RXDLYSRESET);
  buf B_RXELECIDLEMODE0 (RXELECIDLEMODE_IN[0], RXELECIDLEMODE[0]);
  buf B_RXELECIDLEMODE1 (RXELECIDLEMODE_IN[1], RXELECIDLEMODE[1]);
  buf B_RXGEARBOXSLIP (RXGEARBOXSLIP_IN, RXGEARBOXSLIP);
  buf B_RXLPMEN (RXLPMEN_IN, RXLPMEN);
  buf B_RXLPMHFHOLD (RXLPMHFHOLD_IN, RXLPMHFHOLD);
  buf B_RXLPMHFOVRDEN (RXLPMHFOVRDEN_IN, RXLPMHFOVRDEN);
  buf B_RXLPMLFHOLD (RXLPMLFHOLD_IN, RXLPMLFHOLD);
  buf B_RXLPMLFKLOVRDEN (RXLPMLFKLOVRDEN_IN, RXLPMLFKLOVRDEN);
  buf B_RXMCOMMAALIGNEN (RXMCOMMAALIGNEN_IN, RXMCOMMAALIGNEN);
  buf B_RXMONITORSEL0 (RXMONITORSEL_IN[0], RXMONITORSEL[0]);
  buf B_RXMONITORSEL1 (RXMONITORSEL_IN[1], RXMONITORSEL[1]);
  buf B_RXOOBRESET (RXOOBRESET_IN, RXOOBRESET);
  buf B_RXOSHOLD (RXOSHOLD_IN, RXOSHOLD);
  buf B_RXOSOVRDEN (RXOSOVRDEN_IN, RXOSOVRDEN);
  buf B_RXOUTCLKSEL0 (RXOUTCLKSEL_IN[0], RXOUTCLKSEL[0]);
  buf B_RXOUTCLKSEL1 (RXOUTCLKSEL_IN[1], RXOUTCLKSEL[1]);
  buf B_RXOUTCLKSEL2 (RXOUTCLKSEL_IN[2], RXOUTCLKSEL[2]);
  buf B_RXPCOMMAALIGNEN (RXPCOMMAALIGNEN_IN, RXPCOMMAALIGNEN);
  buf B_RXPCSRESET (RXPCSRESET_IN, RXPCSRESET);
  buf B_RXPD0 (RXPD_IN[0], RXPD[0]);
  buf B_RXPD1 (RXPD_IN[1], RXPD[1]);
  buf B_RXPHALIGN (RXPHALIGN_IN, RXPHALIGN);
  buf B_RXPHALIGNEN (RXPHALIGNEN_IN, RXPHALIGNEN);
  buf B_RXPHDLYPD (RXPHDLYPD_IN, RXPHDLYPD);
  buf B_RXPHDLYRESET (RXPHDLYRESET_IN, RXPHDLYRESET);
  buf B_RXPHOVRDEN (RXPHOVRDEN_IN, RXPHOVRDEN);
  buf B_RXPMARESET (RXPMARESET_IN, RXPMARESET);
  buf B_RXPOLARITY (RXPOLARITY_IN, RXPOLARITY);
  buf B_RXPRBSCNTRESET (RXPRBSCNTRESET_IN, RXPRBSCNTRESET);
  buf B_RXPRBSSEL0 (RXPRBSSEL_IN[0], RXPRBSSEL[0]);
  buf B_RXPRBSSEL1 (RXPRBSSEL_IN[1], RXPRBSSEL[1]);
  buf B_RXPRBSSEL2 (RXPRBSSEL_IN[2], RXPRBSSEL[2]);
  buf B_RXQPIEN (RXQPIEN_IN, RXQPIEN);
  buf B_RXRATE0 (RXRATE_IN[0], RXRATE[0]);
  buf B_RXRATE1 (RXRATE_IN[1], RXRATE[1]);
  buf B_RXRATE2 (RXRATE_IN[2], RXRATE[2]);
  buf B_RXSLIDE (RXSLIDE_IN, RXSLIDE);
  buf B_RXSYSCLKSEL0 (RXSYSCLKSEL_IN[0], RXSYSCLKSEL[0]);
  buf B_RXSYSCLKSEL1 (RXSYSCLKSEL_IN[1], RXSYSCLKSEL[1]);
  buf B_RXUSERRDY (RXUSERRDY_IN, RXUSERRDY);
  buf B_RXUSRCLK (RXUSRCLK_IN, RXUSRCLK);
  buf B_RXUSRCLK2 (RXUSRCLK2_IN, RXUSRCLK2);
  buf B_SETERRSTATUS (SETERRSTATUS_IN, SETERRSTATUS);
  buf B_TSTIN0 (TSTIN_IN[0], TSTIN[0]);
  buf B_TSTIN1 (TSTIN_IN[1], TSTIN[1]);
  buf B_TSTIN10 (TSTIN_IN[10], TSTIN[10]);
  buf B_TSTIN11 (TSTIN_IN[11], TSTIN[11]);
  buf B_TSTIN12 (TSTIN_IN[12], TSTIN[12]);
  buf B_TSTIN13 (TSTIN_IN[13], TSTIN[13]);
  buf B_TSTIN14 (TSTIN_IN[14], TSTIN[14]);
  buf B_TSTIN15 (TSTIN_IN[15], TSTIN[15]);
  buf B_TSTIN16 (TSTIN_IN[16], TSTIN[16]);
  buf B_TSTIN17 (TSTIN_IN[17], TSTIN[17]);
  buf B_TSTIN18 (TSTIN_IN[18], TSTIN[18]);
  buf B_TSTIN19 (TSTIN_IN[19], TSTIN[19]);
  buf B_TSTIN2 (TSTIN_IN[2], TSTIN[2]);
  buf B_TSTIN3 (TSTIN_IN[3], TSTIN[3]);
  buf B_TSTIN4 (TSTIN_IN[4], TSTIN[4]);
  buf B_TSTIN5 (TSTIN_IN[5], TSTIN[5]);
  buf B_TSTIN6 (TSTIN_IN[6], TSTIN[6]);
  buf B_TSTIN7 (TSTIN_IN[7], TSTIN[7]);
  buf B_TSTIN8 (TSTIN_IN[8], TSTIN[8]);
  buf B_TSTIN9 (TSTIN_IN[9], TSTIN[9]);
  buf B_TX8B10BBYPASS0 (TX8B10BBYPASS_IN[0], TX8B10BBYPASS[0]);
  buf B_TX8B10BBYPASS1 (TX8B10BBYPASS_IN[1], TX8B10BBYPASS[1]);
  buf B_TX8B10BBYPASS2 (TX8B10BBYPASS_IN[2], TX8B10BBYPASS[2]);
  buf B_TX8B10BBYPASS3 (TX8B10BBYPASS_IN[3], TX8B10BBYPASS[3]);
  buf B_TX8B10BBYPASS4 (TX8B10BBYPASS_IN[4], TX8B10BBYPASS[4]);
  buf B_TX8B10BBYPASS5 (TX8B10BBYPASS_IN[5], TX8B10BBYPASS[5]);
  buf B_TX8B10BBYPASS6 (TX8B10BBYPASS_IN[6], TX8B10BBYPASS[6]);
  buf B_TX8B10BBYPASS7 (TX8B10BBYPASS_IN[7], TX8B10BBYPASS[7]);
  buf B_TX8B10BEN (TX8B10BEN_IN, TX8B10BEN);
  buf B_TXBUFDIFFCTRL0 (TXBUFDIFFCTRL_IN[0], TXBUFDIFFCTRL[0]);
  buf B_TXBUFDIFFCTRL1 (TXBUFDIFFCTRL_IN[1], TXBUFDIFFCTRL[1]);
  buf B_TXBUFDIFFCTRL2 (TXBUFDIFFCTRL_IN[2], TXBUFDIFFCTRL[2]);
  buf B_TXCHARDISPMODE0 (TXCHARDISPMODE_IN[0], TXCHARDISPMODE[0]);
  buf B_TXCHARDISPMODE1 (TXCHARDISPMODE_IN[1], TXCHARDISPMODE[1]);
  buf B_TXCHARDISPMODE2 (TXCHARDISPMODE_IN[2], TXCHARDISPMODE[2]);
  buf B_TXCHARDISPMODE3 (TXCHARDISPMODE_IN[3], TXCHARDISPMODE[3]);
  buf B_TXCHARDISPMODE4 (TXCHARDISPMODE_IN[4], TXCHARDISPMODE[4]);
  buf B_TXCHARDISPMODE5 (TXCHARDISPMODE_IN[5], TXCHARDISPMODE[5]);
  buf B_TXCHARDISPMODE6 (TXCHARDISPMODE_IN[6], TXCHARDISPMODE[6]);
  buf B_TXCHARDISPMODE7 (TXCHARDISPMODE_IN[7], TXCHARDISPMODE[7]);
  buf B_TXCHARDISPVAL0 (TXCHARDISPVAL_IN[0], TXCHARDISPVAL[0]);
  buf B_TXCHARDISPVAL1 (TXCHARDISPVAL_IN[1], TXCHARDISPVAL[1]);
  buf B_TXCHARDISPVAL2 (TXCHARDISPVAL_IN[2], TXCHARDISPVAL[2]);
  buf B_TXCHARDISPVAL3 (TXCHARDISPVAL_IN[3], TXCHARDISPVAL[3]);
  buf B_TXCHARDISPVAL4 (TXCHARDISPVAL_IN[4], TXCHARDISPVAL[4]);
  buf B_TXCHARDISPVAL5 (TXCHARDISPVAL_IN[5], TXCHARDISPVAL[5]);
  buf B_TXCHARDISPVAL6 (TXCHARDISPVAL_IN[6], TXCHARDISPVAL[6]);
  buf B_TXCHARDISPVAL7 (TXCHARDISPVAL_IN[7], TXCHARDISPVAL[7]);
  buf B_TXCHARISK0 (TXCHARISK_IN[0], TXCHARISK[0]);
  buf B_TXCHARISK1 (TXCHARISK_IN[1], TXCHARISK[1]);
  buf B_TXCHARISK2 (TXCHARISK_IN[2], TXCHARISK[2]);
  buf B_TXCHARISK3 (TXCHARISK_IN[3], TXCHARISK[3]);
  buf B_TXCHARISK4 (TXCHARISK_IN[4], TXCHARISK[4]);
  buf B_TXCHARISK5 (TXCHARISK_IN[5], TXCHARISK[5]);
  buf B_TXCHARISK6 (TXCHARISK_IN[6], TXCHARISK[6]);
  buf B_TXCHARISK7 (TXCHARISK_IN[7], TXCHARISK[7]);
  buf B_TXCOMINIT (TXCOMINIT_IN, TXCOMINIT);
  buf B_TXCOMSAS (TXCOMSAS_IN, TXCOMSAS);
  buf B_TXCOMWAKE (TXCOMWAKE_IN, TXCOMWAKE);
  buf B_TXDATA0 (TXDATA_IN[0], TXDATA[0]);
  buf B_TXDATA1 (TXDATA_IN[1], TXDATA[1]);
  buf B_TXDATA10 (TXDATA_IN[10], TXDATA[10]);
  buf B_TXDATA11 (TXDATA_IN[11], TXDATA[11]);
  buf B_TXDATA12 (TXDATA_IN[12], TXDATA[12]);
  buf B_TXDATA13 (TXDATA_IN[13], TXDATA[13]);
  buf B_TXDATA14 (TXDATA_IN[14], TXDATA[14]);
  buf B_TXDATA15 (TXDATA_IN[15], TXDATA[15]);
  buf B_TXDATA16 (TXDATA_IN[16], TXDATA[16]);
  buf B_TXDATA17 (TXDATA_IN[17], TXDATA[17]);
  buf B_TXDATA18 (TXDATA_IN[18], TXDATA[18]);
  buf B_TXDATA19 (TXDATA_IN[19], TXDATA[19]);
  buf B_TXDATA2 (TXDATA_IN[2], TXDATA[2]);
  buf B_TXDATA20 (TXDATA_IN[20], TXDATA[20]);
  buf B_TXDATA21 (TXDATA_IN[21], TXDATA[21]);
  buf B_TXDATA22 (TXDATA_IN[22], TXDATA[22]);
  buf B_TXDATA23 (TXDATA_IN[23], TXDATA[23]);
  buf B_TXDATA24 (TXDATA_IN[24], TXDATA[24]);
  buf B_TXDATA25 (TXDATA_IN[25], TXDATA[25]);
  buf B_TXDATA26 (TXDATA_IN[26], TXDATA[26]);
  buf B_TXDATA27 (TXDATA_IN[27], TXDATA[27]);
  buf B_TXDATA28 (TXDATA_IN[28], TXDATA[28]);
  buf B_TXDATA29 (TXDATA_IN[29], TXDATA[29]);
  buf B_TXDATA3 (TXDATA_IN[3], TXDATA[3]);
  buf B_TXDATA30 (TXDATA_IN[30], TXDATA[30]);
  buf B_TXDATA31 (TXDATA_IN[31], TXDATA[31]);
  buf B_TXDATA32 (TXDATA_IN[32], TXDATA[32]);
  buf B_TXDATA33 (TXDATA_IN[33], TXDATA[33]);
  buf B_TXDATA34 (TXDATA_IN[34], TXDATA[34]);
  buf B_TXDATA35 (TXDATA_IN[35], TXDATA[35]);
  buf B_TXDATA36 (TXDATA_IN[36], TXDATA[36]);
  buf B_TXDATA37 (TXDATA_IN[37], TXDATA[37]);
  buf B_TXDATA38 (TXDATA_IN[38], TXDATA[38]);
  buf B_TXDATA39 (TXDATA_IN[39], TXDATA[39]);
  buf B_TXDATA4 (TXDATA_IN[4], TXDATA[4]);
  buf B_TXDATA40 (TXDATA_IN[40], TXDATA[40]);
  buf B_TXDATA41 (TXDATA_IN[41], TXDATA[41]);
  buf B_TXDATA42 (TXDATA_IN[42], TXDATA[42]);
  buf B_TXDATA43 (TXDATA_IN[43], TXDATA[43]);
  buf B_TXDATA44 (TXDATA_IN[44], TXDATA[44]);
  buf B_TXDATA45 (TXDATA_IN[45], TXDATA[45]);
  buf B_TXDATA46 (TXDATA_IN[46], TXDATA[46]);
  buf B_TXDATA47 (TXDATA_IN[47], TXDATA[47]);
  buf B_TXDATA48 (TXDATA_IN[48], TXDATA[48]);
  buf B_TXDATA49 (TXDATA_IN[49], TXDATA[49]);
  buf B_TXDATA5 (TXDATA_IN[5], TXDATA[5]);
  buf B_TXDATA50 (TXDATA_IN[50], TXDATA[50]);
  buf B_TXDATA51 (TXDATA_IN[51], TXDATA[51]);
  buf B_TXDATA52 (TXDATA_IN[52], TXDATA[52]);
  buf B_TXDATA53 (TXDATA_IN[53], TXDATA[53]);
  buf B_TXDATA54 (TXDATA_IN[54], TXDATA[54]);
  buf B_TXDATA55 (TXDATA_IN[55], TXDATA[55]);
  buf B_TXDATA56 (TXDATA_IN[56], TXDATA[56]);
  buf B_TXDATA57 (TXDATA_IN[57], TXDATA[57]);
  buf B_TXDATA58 (TXDATA_IN[58], TXDATA[58]);
  buf B_TXDATA59 (TXDATA_IN[59], TXDATA[59]);
  buf B_TXDATA6 (TXDATA_IN[6], TXDATA[6]);
  buf B_TXDATA60 (TXDATA_IN[60], TXDATA[60]);
  buf B_TXDATA61 (TXDATA_IN[61], TXDATA[61]);
  buf B_TXDATA62 (TXDATA_IN[62], TXDATA[62]);
  buf B_TXDATA63 (TXDATA_IN[63], TXDATA[63]);
  buf B_TXDATA7 (TXDATA_IN[7], TXDATA[7]);
  buf B_TXDATA8 (TXDATA_IN[8], TXDATA[8]);
  buf B_TXDATA9 (TXDATA_IN[9], TXDATA[9]);
  buf B_TXDEEMPH (TXDEEMPH_IN, TXDEEMPH);
  buf B_TXDETECTRX (TXDETECTRX_IN, TXDETECTRX);
  buf B_TXDIFFCTRL0 (TXDIFFCTRL_IN[0], TXDIFFCTRL[0]);
  buf B_TXDIFFCTRL1 (TXDIFFCTRL_IN[1], TXDIFFCTRL[1]);
  buf B_TXDIFFCTRL2 (TXDIFFCTRL_IN[2], TXDIFFCTRL[2]);
  buf B_TXDIFFCTRL3 (TXDIFFCTRL_IN[3], TXDIFFCTRL[3]);
  buf B_TXDIFFPD (TXDIFFPD_IN, TXDIFFPD);
  buf B_TXDLYBYPASS (TXDLYBYPASS_IN, TXDLYBYPASS);
  buf B_TXDLYEN (TXDLYEN_IN, TXDLYEN);
  buf B_TXDLYHOLD (TXDLYHOLD_IN, TXDLYHOLD);
  buf B_TXDLYOVRDEN (TXDLYOVRDEN_IN, TXDLYOVRDEN);
  buf B_TXDLYSRESET (TXDLYSRESET_IN, TXDLYSRESET);
  buf B_TXDLYUPDOWN (TXDLYUPDOWN_IN, TXDLYUPDOWN);
  buf B_TXELECIDLE (TXELECIDLE_IN, TXELECIDLE);
  buf B_TXHEADER0 (TXHEADER_IN[0], TXHEADER[0]);
  buf B_TXHEADER1 (TXHEADER_IN[1], TXHEADER[1]);
  buf B_TXHEADER2 (TXHEADER_IN[2], TXHEADER[2]);
  buf B_TXINHIBIT (TXINHIBIT_IN, TXINHIBIT);
  buf B_TXMAINCURSOR0 (TXMAINCURSOR_IN[0], TXMAINCURSOR[0]);
  buf B_TXMAINCURSOR1 (TXMAINCURSOR_IN[1], TXMAINCURSOR[1]);
  buf B_TXMAINCURSOR2 (TXMAINCURSOR_IN[2], TXMAINCURSOR[2]);
  buf B_TXMAINCURSOR3 (TXMAINCURSOR_IN[3], TXMAINCURSOR[3]);
  buf B_TXMAINCURSOR4 (TXMAINCURSOR_IN[4], TXMAINCURSOR[4]);
  buf B_TXMAINCURSOR5 (TXMAINCURSOR_IN[5], TXMAINCURSOR[5]);
  buf B_TXMAINCURSOR6 (TXMAINCURSOR_IN[6], TXMAINCURSOR[6]);
  buf B_TXMARGIN0 (TXMARGIN_IN[0], TXMARGIN[0]);
  buf B_TXMARGIN1 (TXMARGIN_IN[1], TXMARGIN[1]);
  buf B_TXMARGIN2 (TXMARGIN_IN[2], TXMARGIN[2]);
  buf B_TXOUTCLKSEL0 (TXOUTCLKSEL_IN[0], TXOUTCLKSEL[0]);
  buf B_TXOUTCLKSEL1 (TXOUTCLKSEL_IN[1], TXOUTCLKSEL[1]);
  buf B_TXOUTCLKSEL2 (TXOUTCLKSEL_IN[2], TXOUTCLKSEL[2]);
  buf B_TXPCSRESET (TXPCSRESET_IN, TXPCSRESET);
  buf B_TXPD0 (TXPD_IN[0], TXPD[0]);
  buf B_TXPD1 (TXPD_IN[1], TXPD[1]);
  buf B_TXPDELECIDLEMODE (TXPDELECIDLEMODE_IN, TXPDELECIDLEMODE);
  buf B_TXPHALIGN (TXPHALIGN_IN, TXPHALIGN);
  buf B_TXPHALIGNEN (TXPHALIGNEN_IN, TXPHALIGNEN);
  buf B_TXPHDLYPD (TXPHDLYPD_IN, TXPHDLYPD);
  buf B_TXPHDLYRESET (TXPHDLYRESET_IN, TXPHDLYRESET);
  buf B_TXPHDLYTSTCLK (TXPHDLYTSTCLK_IN, TXPHDLYTSTCLK);
  buf B_TXPHINIT (TXPHINIT_IN, TXPHINIT);
  buf B_TXPHOVRDEN (TXPHOVRDEN_IN, TXPHOVRDEN);
  buf B_TXPISOPD (TXPISOPD_IN, TXPISOPD);
  buf B_TXPMARESET (TXPMARESET_IN, TXPMARESET);
  buf B_TXPOLARITY (TXPOLARITY_IN, TXPOLARITY);
  buf B_TXPOSTCURSOR0 (TXPOSTCURSOR_IN[0], TXPOSTCURSOR[0]);
  buf B_TXPOSTCURSOR1 (TXPOSTCURSOR_IN[1], TXPOSTCURSOR[1]);
  buf B_TXPOSTCURSOR2 (TXPOSTCURSOR_IN[2], TXPOSTCURSOR[2]);
  buf B_TXPOSTCURSOR3 (TXPOSTCURSOR_IN[3], TXPOSTCURSOR[3]);
  buf B_TXPOSTCURSOR4 (TXPOSTCURSOR_IN[4], TXPOSTCURSOR[4]);
  buf B_TXPOSTCURSORINV (TXPOSTCURSORINV_IN, TXPOSTCURSORINV);
  buf B_TXPRBSFORCEERR (TXPRBSFORCEERR_IN, TXPRBSFORCEERR);
  buf B_TXPRBSSEL0 (TXPRBSSEL_IN[0], TXPRBSSEL[0]);
  buf B_TXPRBSSEL1 (TXPRBSSEL_IN[1], TXPRBSSEL[1]);
  buf B_TXPRBSSEL2 (TXPRBSSEL_IN[2], TXPRBSSEL[2]);
  buf B_TXPRECURSOR0 (TXPRECURSOR_IN[0], TXPRECURSOR[0]);
  buf B_TXPRECURSOR1 (TXPRECURSOR_IN[1], TXPRECURSOR[1]);
  buf B_TXPRECURSOR2 (TXPRECURSOR_IN[2], TXPRECURSOR[2]);
  buf B_TXPRECURSOR3 (TXPRECURSOR_IN[3], TXPRECURSOR[3]);
  buf B_TXPRECURSOR4 (TXPRECURSOR_IN[4], TXPRECURSOR[4]);
  buf B_TXPRECURSORINV (TXPRECURSORINV_IN, TXPRECURSORINV);
  buf B_TXQPIBIASEN (TXQPIBIASEN_IN, TXQPIBIASEN);
  buf B_TXQPISTRONGPDOWN (TXQPISTRONGPDOWN_IN, TXQPISTRONGPDOWN);
  buf B_TXQPIWEAKPUP (TXQPIWEAKPUP_IN, TXQPIWEAKPUP);
  buf B_TXRATE0 (TXRATE_IN[0], TXRATE[0]);
  buf B_TXRATE1 (TXRATE_IN[1], TXRATE[1]);
  buf B_TXRATE2 (TXRATE_IN[2], TXRATE[2]);
  buf B_TXSEQUENCE0 (TXSEQUENCE_IN[0], TXSEQUENCE[0]);
  buf B_TXSEQUENCE1 (TXSEQUENCE_IN[1], TXSEQUENCE[1]);
  buf B_TXSEQUENCE2 (TXSEQUENCE_IN[2], TXSEQUENCE[2]);
  buf B_TXSEQUENCE3 (TXSEQUENCE_IN[3], TXSEQUENCE[3]);
  buf B_TXSEQUENCE4 (TXSEQUENCE_IN[4], TXSEQUENCE[4]);
  buf B_TXSEQUENCE5 (TXSEQUENCE_IN[5], TXSEQUENCE[5]);
  buf B_TXSEQUENCE6 (TXSEQUENCE_IN[6], TXSEQUENCE[6]);
  buf B_TXSTARTSEQ (TXSTARTSEQ_IN, TXSTARTSEQ);
  buf B_TXSWING (TXSWING_IN, TXSWING);
  buf B_TXSYSCLKSEL0 (TXSYSCLKSEL_IN[0], TXSYSCLKSEL[0]);
  buf B_TXSYSCLKSEL1 (TXSYSCLKSEL_IN[1], TXSYSCLKSEL[1]);
  buf B_TXUSERRDY (TXUSERRDY_IN, TXUSERRDY);
  buf B_TXUSRCLK (TXUSRCLK_IN, TXUSRCLK);
  buf B_TXUSRCLK2 (TXUSRCLK2_IN, TXUSRCLK2);

  wire [15:0] delay_DRPDO;
  wire [15:0] delay_PCSRSVDOUT;
  wire [1:0] delay_RXCLKCORCNT;
  wire [1:0] delay_TXBUFSTATUS;
  wire [2:0] delay_RXBUFSTATUS;
  wire [2:0] delay_RXHEADER;
  wire [2:0] delay_RXSTATUS;
  wire [4:0] delay_RXCHBONDO;
  wire [4:0] delay_RXPHMONITOR;
  wire [4:0] delay_RXPHSLIPMONITOR;
  wire [63:0] delay_RXDATA;
  wire [6:0] delay_RXMONITOROUT;
  wire [7:0] delay_DMONITOROUT;
  wire [7:0] delay_RXCHARISCOMMA;
  wire [7:0] delay_RXCHARISK;
  wire [7:0] delay_RXDISPERR;
  wire [7:0] delay_RXNOTINTABLE;
  wire [9:0] delay_TSTOUT;
  wire delay_CPLLFBCLKLOST;
  wire delay_CPLLLOCK;
  wire delay_CPLLREFCLKLOST;
  wire delay_DRPRDY;
  wire delay_EYESCANDATAERROR;
  wire delay_GTREFCLKMONITOR;
  wire delay_GTXTXN;
  wire delay_GTXTXP;
  wire delay_PHYSTATUS;
  wire delay_RXBYTEISALIGNED;
  wire delay_RXBYTEREALIGN;
  wire delay_RXCDRLOCK;
  wire delay_RXCHANBONDSEQ;
  wire delay_RXCHANISALIGNED;
  wire delay_RXCHANREALIGN;
  wire delay_RXCOMINITDET;
  wire delay_RXCOMMADET;
  wire delay_RXCOMSASDET;
  wire delay_RXCOMWAKEDET;
  wire delay_RXDATAVALID;
  wire delay_RXDLYSRESETDONE;
  wire delay_RXELECIDLE;
  wire delay_RXHEADERVALID;
  wire delay_RXOUTCLK;
  wire delay_RXOUTCLKFABRIC;
  wire delay_RXOUTCLKPCS;
  wire delay_RXPHALIGNDONE;
  wire delay_RXPRBSERR;
  wire delay_RXQPISENN;
  wire delay_RXQPISENP;
  wire delay_RXRATEDONE;
  wire delay_RXRESETDONE;
  wire delay_RXSTARTOFSEQ;
  wire delay_RXVALID;
  wire delay_TXCOMFINISH;
  wire delay_TXDLYSRESETDONE;
  wire delay_TXGEARBOXREADY;
  wire delay_TXOUTCLK;
  wire delay_TXOUTCLKFABRIC;
  wire delay_TXOUTCLKPCS;
  wire delay_TXPHALIGNDONE;
  wire delay_TXPHINITDONE;
  wire delay_TXQPISENN;
  wire delay_TXQPISENP;
  wire delay_TXRATEDONE;
  wire delay_TXRESETDONE;

  wire [15:0] delay_DRPDI;
  wire [15:0] delay_GTRSVD;
  wire [15:0] delay_PCSRSVDIN;
  wire [19:0] delay_TSTIN;
  wire [1:0] delay_RXELECIDLEMODE;
  wire [1:0] delay_RXMONITORSEL;
  wire [1:0] delay_RXPD;
  wire [1:0] delay_RXSYSCLKSEL;
  wire [1:0] delay_TXPD;
  wire [1:0] delay_TXSYSCLKSEL;
  wire [2:0] delay_CPLLREFCLKSEL;
  wire [2:0] delay_LOOPBACK;
  wire [2:0] delay_RXCHBONDLEVEL;
  wire [2:0] delay_RXOUTCLKSEL;
  wire [2:0] delay_RXPRBSSEL;
  wire [2:0] delay_RXRATE;
  wire [2:0] delay_TXBUFDIFFCTRL;
  wire [2:0] delay_TXHEADER;
  wire [2:0] delay_TXMARGIN;
  wire [2:0] delay_TXOUTCLKSEL;
  wire [2:0] delay_TXPRBSSEL;
  wire [2:0] delay_TXRATE;
  wire [3:0] delay_CLKRSVD;
  wire [3:0] delay_TXDIFFCTRL;
  wire [4:0] delay_PCSRSVDIN2;
  wire [4:0] delay_PMARSVDIN2;
  wire [4:0] delay_PMARSVDIN;
  wire [4:0] delay_RXCHBONDI;
  wire [4:0] delay_TXPOSTCURSOR;
  wire [4:0] delay_TXPRECURSOR;
  wire [63:0] delay_TXDATA;
  wire [6:0] delay_TXMAINCURSOR;
  wire [6:0] delay_TXSEQUENCE;
  wire [7:0] delay_TX8B10BBYPASS;
  wire [7:0] delay_TXCHARDISPMODE;
  wire [7:0] delay_TXCHARDISPVAL;
  wire [7:0] delay_TXCHARISK;
  wire [8:0] delay_DRPADDR;
  wire delay_CFGRESET;
  wire delay_CPLLLOCKDETCLK;
  wire delay_CPLLLOCKEN;
  wire delay_CPLLPD;
  wire delay_CPLLRESET;
  wire delay_DRPCLK;
  wire delay_DRPEN;
  wire delay_DRPWE;
  wire delay_EYESCANMODE;
  wire delay_EYESCANRESET;
  wire delay_EYESCANTRIGGER;
  wire delay_GTGREFCLK;
  wire delay_GTNORTHREFCLK0;
  wire delay_GTNORTHREFCLK1;
  wire delay_GTREFCLK0;
  wire delay_GTREFCLK1;
  wire delay_GTRESETSEL;
  wire delay_GTRXRESET;
  wire delay_GTSOUTHREFCLK0;
  wire delay_GTSOUTHREFCLK1;
  wire delay_GTTXRESET;
  wire delay_GTXRXN;
  wire delay_GTXRXP;
  wire delay_QPLLCLK;
  wire delay_QPLLREFCLK;
  wire delay_RESETOVRD;
  wire delay_RX8B10BEN;
  wire delay_RXBUFRESET;
  wire delay_RXCDRFREQRESET;
  wire delay_RXCDRHOLD;
  wire delay_RXCDROVRDEN;
  wire delay_RXCDRRESET;
  wire delay_RXCDRRESETRSV;
  wire delay_RXCHBONDEN;
  wire delay_RXCHBONDMASTER;
  wire delay_RXCHBONDSLAVE;
  wire delay_RXCOMMADETEN;
  wire delay_RXDDIEN;
  wire delay_RXDFEAGCHOLD;
  wire delay_RXDFEAGCOVRDEN;
  wire delay_RXDFECM1EN;
  wire delay_RXDFELFHOLD;
  wire delay_RXDFELFOVRDEN;
  wire delay_RXDFELPMRESET;
  wire delay_RXDFETAP2HOLD;
  wire delay_RXDFETAP2OVRDEN;
  wire delay_RXDFETAP3HOLD;
  wire delay_RXDFETAP3OVRDEN;
  wire delay_RXDFETAP4HOLD;
  wire delay_RXDFETAP4OVRDEN;
  wire delay_RXDFETAP5HOLD;
  wire delay_RXDFETAP5OVRDEN;
  wire delay_RXDFEUTHOLD;
  wire delay_RXDFEUTOVRDEN;
  wire delay_RXDFEVPHOLD;
  wire delay_RXDFEVPOVRDEN;
  wire delay_RXDFEVSEN;
  wire delay_RXDFEXYDEN;
  wire delay_RXDFEXYDHOLD;
  wire delay_RXDFEXYDOVRDEN;
  wire delay_RXDLYBYPASS;
  wire delay_RXDLYEN;
  wire delay_RXDLYOVRDEN;
  wire delay_RXDLYSRESET;
  wire delay_RXGEARBOXSLIP;
  wire delay_RXLPMEN;
  wire delay_RXLPMHFHOLD;
  wire delay_RXLPMHFOVRDEN;
  wire delay_RXLPMLFHOLD;
  wire delay_RXLPMLFKLOVRDEN;
  wire delay_RXMCOMMAALIGNEN;
  wire delay_RXOOBRESET;
  wire delay_RXOSHOLD;
  wire delay_RXOSOVRDEN;
  wire delay_RXPCOMMAALIGNEN;
  wire delay_RXPCSRESET;
  wire delay_RXPHALIGN;
  wire delay_RXPHALIGNEN;
  wire delay_RXPHDLYPD;
  wire delay_RXPHDLYRESET;
  wire delay_RXPHOVRDEN;
  wire delay_RXPMARESET;
  wire delay_RXPOLARITY;
  wire delay_RXPRBSCNTRESET;
  wire delay_RXQPIEN;
  wire delay_RXSLIDE;
  wire delay_RXUSERRDY;
  wire delay_RXUSRCLK2;
  wire delay_RXUSRCLK;
  wire delay_SETERRSTATUS;
  wire delay_TX8B10BEN;
  wire delay_TXCOMINIT;
  wire delay_TXCOMSAS;
  wire delay_TXCOMWAKE;
  wire delay_TXDEEMPH;
  wire delay_TXDETECTRX;
  wire delay_TXDIFFPD;
  wire delay_TXDLYBYPASS;
  wire delay_TXDLYEN;
  wire delay_TXDLYHOLD;
  wire delay_TXDLYOVRDEN;
  wire delay_TXDLYSRESET;
  wire delay_TXDLYUPDOWN;
  wire delay_TXELECIDLE;
  wire delay_TXINHIBIT;
  wire delay_TXPCSRESET;
  wire delay_TXPDELECIDLEMODE;
  wire delay_TXPHALIGN;
  wire delay_TXPHALIGNEN;
  wire delay_TXPHDLYPD;
  wire delay_TXPHDLYRESET;
  wire delay_TXPHDLYTSTCLK;
  wire delay_TXPHINIT;
  wire delay_TXPHOVRDEN;
  wire delay_TXPISOPD;
  wire delay_TXPMARESET;
  wire delay_TXPOLARITY;
  wire delay_TXPOSTCURSORINV;
  wire delay_TXPRBSFORCEERR;
  wire delay_TXPRECURSORINV;
  wire delay_TXQPIBIASEN;
  wire delay_TXQPISTRONGPDOWN;
  wire delay_TXQPIWEAKPUP;
  wire delay_TXSTARTSEQ;
  wire delay_TXSWING;
  wire delay_TXUSERRDY;
  wire delay_TXUSRCLK2;
  wire delay_TXUSRCLK;

  assign #(OUTCLK_DELAY) GTREFCLKMONITOR_OUT = delay_GTREFCLKMONITOR;
  assign #(OUTCLK_DELAY) RXOUTCLK_OUT = delay_RXOUTCLK;
  assign #(OUTCLK_DELAY) TXOUTCLK_OUT = delay_TXOUTCLK;

  assign #(out_delay) CPLLFBCLKLOST_OUT = delay_CPLLFBCLKLOST;
  assign #(out_delay) CPLLLOCK_OUT = delay_CPLLLOCK;
  assign #(out_delay) CPLLREFCLKLOST_OUT = delay_CPLLREFCLKLOST;
  assign #(out_delay) DMONITOROUT_OUT = delay_DMONITOROUT;
  assign #(out_delay) DRPDO_OUT = delay_DRPDO;
  assign #(out_delay) DRPRDY_OUT = delay_DRPRDY;
  assign #(out_delay) EYESCANDATAERROR_OUT = delay_EYESCANDATAERROR;
  assign #(out_delay) GTXTXN_OUT = delay_GTXTXN;
  assign #(out_delay) GTXTXP_OUT = delay_GTXTXP;
  assign #(out_delay) PCSRSVDOUT_OUT = delay_PCSRSVDOUT;
  assign #(out_delay) PHYSTATUS_OUT = delay_PHYSTATUS;
  assign #(out_delay) RXBUFSTATUS_OUT = delay_RXBUFSTATUS;
  assign #(out_delay) RXBYTEISALIGNED_OUT = delay_RXBYTEISALIGNED;
  assign #(out_delay) RXBYTEREALIGN_OUT = delay_RXBYTEREALIGN;
  assign #(out_delay) RXCDRLOCK_OUT = delay_RXCDRLOCK;
  assign #(out_delay) RXCHANBONDSEQ_OUT = delay_RXCHANBONDSEQ;
  assign #(out_delay) RXCHANISALIGNED_OUT = delay_RXCHANISALIGNED;
  assign #(out_delay) RXCHANREALIGN_OUT = delay_RXCHANREALIGN;
  assign #(out_delay) RXCHARISCOMMA_OUT = delay_RXCHARISCOMMA;
  assign #(out_delay) RXCHARISK_OUT = delay_RXCHARISK;
  assign #(out_delay) RXCHBONDO_OUT = delay_RXCHBONDO;
  assign #(out_delay) RXCLKCORCNT_OUT = delay_RXCLKCORCNT;
  assign #(out_delay) RXCOMINITDET_OUT = delay_RXCOMINITDET;
  assign #(out_delay) RXCOMMADET_OUT = delay_RXCOMMADET;
  assign #(out_delay) RXCOMSASDET_OUT = delay_RXCOMSASDET;
  assign #(out_delay) RXCOMWAKEDET_OUT = delay_RXCOMWAKEDET;
  assign #(out_delay) RXDATAVALID_OUT = delay_RXDATAVALID;
  assign #(out_delay) RXDATA_OUT = delay_RXDATA;
  assign #(out_delay) RXDISPERR_OUT = delay_RXDISPERR;
  assign #(out_delay) RXDLYSRESETDONE_OUT = delay_RXDLYSRESETDONE;
  assign #(out_delay) RXELECIDLE_OUT = delay_RXELECIDLE;
  assign #(out_delay) RXHEADERVALID_OUT = delay_RXHEADERVALID;
  assign #(out_delay) RXHEADER_OUT = delay_RXHEADER;
  assign #(out_delay) RXMONITOROUT_OUT = delay_RXMONITOROUT;
  assign #(out_delay) RXNOTINTABLE_OUT = delay_RXNOTINTABLE;
  assign #(out_delay) RXOUTCLKFABRIC_OUT = delay_RXOUTCLKFABRIC;
  assign #(out_delay) RXOUTCLKPCS_OUT = delay_RXOUTCLKPCS;
  assign #(out_delay) RXPHALIGNDONE_OUT = delay_RXPHALIGNDONE;
  assign #(out_delay) RXPHMONITOR_OUT = delay_RXPHMONITOR;
  assign #(out_delay) RXPHSLIPMONITOR_OUT = delay_RXPHSLIPMONITOR;
  assign #(out_delay) RXPRBSERR_OUT = delay_RXPRBSERR;
  assign #(out_delay) RXQPISENN_OUT = delay_RXQPISENN;
  assign #(out_delay) RXQPISENP_OUT = delay_RXQPISENP;
  assign #(out_delay) RXRATEDONE_OUT = delay_RXRATEDONE;
  assign #(out_delay) RXRESETDONE_OUT = delay_RXRESETDONE;
  assign #(out_delay) RXSTARTOFSEQ_OUT = delay_RXSTARTOFSEQ;
  assign #(out_delay) RXSTATUS_OUT = delay_RXSTATUS;
  assign #(out_delay) RXVALID_OUT = delay_RXVALID;
  assign #(out_delay) TSTOUT_OUT = delay_TSTOUT;
  assign #(out_delay) TXBUFSTATUS_OUT = delay_TXBUFSTATUS;
  assign #(out_delay) TXCOMFINISH_OUT = delay_TXCOMFINISH;
  assign #(out_delay) TXDLYSRESETDONE_OUT = delay_TXDLYSRESETDONE;
  assign #(out_delay) TXGEARBOXREADY_OUT = delay_TXGEARBOXREADY;
  assign #(out_delay) TXOUTCLKFABRIC_OUT = delay_TXOUTCLKFABRIC;
  assign #(out_delay) TXOUTCLKPCS_OUT = delay_TXOUTCLKPCS;
  assign #(out_delay) TXPHALIGNDONE_OUT = delay_TXPHALIGNDONE;
  assign #(out_delay) TXPHINITDONE_OUT = delay_TXPHINITDONE;
  assign #(out_delay) TXQPISENN_OUT = delay_TXQPISENN;
  assign #(out_delay) TXQPISENP_OUT = delay_TXQPISENP;
  assign #(out_delay) TXRATEDONE_OUT = delay_TXRATEDONE;
  assign #(out_delay) TXRESETDONE_OUT = delay_TXRESETDONE;

  assign #(INCLK_DELAY) CPLLLOCKDETCLK_INDELAY = CPLLLOCKDETCLK_IN;
  assign #(INCLK_DELAY) DRPCLK_INDELAY = DRPCLK_IN;
  assign #(INCLK_DELAY) GTGREFCLK_INDELAY = GTGREFCLK_IN;
  assign #(INCLK_DELAY) GTNORTHREFCLK0_INDELAY = GTNORTHREFCLK0_IN;
  assign #(INCLK_DELAY) GTNORTHREFCLK1_INDELAY = GTNORTHREFCLK1_IN;
  assign #(INCLK_DELAY) GTREFCLK0_INDELAY = GTREFCLK0_IN;
  assign #(INCLK_DELAY) GTREFCLK1_INDELAY = GTREFCLK1_IN;
  assign #(INCLK_DELAY) GTSOUTHREFCLK0_INDELAY = GTSOUTHREFCLK0_IN;
  assign #(INCLK_DELAY) GTSOUTHREFCLK1_INDELAY = GTSOUTHREFCLK1_IN;
  assign #(INCLK_DELAY) QPLLCLK_INDELAY = QPLLCLK_IN;
  assign #(INCLK_DELAY) RXUSRCLK2_INDELAY = RXUSRCLK2_IN;
  assign #(INCLK_DELAY) RXUSRCLK_INDELAY = RXUSRCLK_IN;
  assign #(INCLK_DELAY) TXPHDLYTSTCLK_INDELAY = TXPHDLYTSTCLK_IN;
  assign #(INCLK_DELAY) TXUSRCLK2_INDELAY = TXUSRCLK2_IN;
  assign #(INCLK_DELAY) TXUSRCLK_INDELAY = TXUSRCLK_IN;

  assign #(in_delay) CFGRESET_INDELAY = CFGRESET_IN;
  assign #(in_delay) CLKRSVD_INDELAY = CLKRSVD_IN;
  assign #(in_delay) CPLLLOCKEN_INDELAY = CPLLLOCKEN_IN;
  assign #(in_delay) CPLLPD_INDELAY = CPLLPD_IN;
  assign #(in_delay) CPLLREFCLKSEL_INDELAY = CPLLREFCLKSEL_IN;
  assign #(in_delay) CPLLRESET_INDELAY = CPLLRESET_IN;
  assign #(in_delay) DRPADDR_INDELAY = DRPADDR_IN;
  assign #(in_delay) DRPDI_INDELAY = DRPDI_IN;
  assign #(in_delay) DRPEN_INDELAY = DRPEN_IN;
  assign #(in_delay) DRPWE_INDELAY = DRPWE_IN;
  assign #(in_delay) EYESCANMODE_INDELAY = EYESCANMODE_IN;
  assign #(in_delay) EYESCANRESET_INDELAY = EYESCANRESET_IN;
  assign #(in_delay) EYESCANTRIGGER_INDELAY = EYESCANTRIGGER_IN;
  assign #(in_delay) GTRESETSEL_INDELAY = GTRESETSEL_IN;
  assign #(in_delay) GTRSVD_INDELAY = GTRSVD_IN;
  assign #(in_delay) GTRXRESET_INDELAY = GTRXRESET_IN;
  assign #(in_delay) GTTXRESET_INDELAY = GTTXRESET_IN;
  assign #(in_delay) GTXRXN_INDELAY = GTXRXN_IN;
  assign #(in_delay) GTXRXP_INDELAY = GTXRXP_IN;
  assign #(in_delay) LOOPBACK_INDELAY = LOOPBACK_IN;
  assign #(in_delay) PCSRSVDIN2_INDELAY = PCSRSVDIN2_IN;
  assign #(in_delay) PCSRSVDIN_INDELAY = PCSRSVDIN_IN;
  assign #(in_delay) PMARSVDIN2_INDELAY = PMARSVDIN2_IN;
  assign #(in_delay) PMARSVDIN_INDELAY = PMARSVDIN_IN;
  assign #(in_delay) QPLLREFCLK_INDELAY = QPLLREFCLK_IN;
  assign #(in_delay) RESETOVRD_INDELAY = RESETOVRD_IN;
  assign #(in_delay) RX8B10BEN_INDELAY = RX8B10BEN_IN;
  assign #(in_delay) RXBUFRESET_INDELAY = RXBUFRESET_IN;
  assign #(in_delay) RXCDRFREQRESET_INDELAY = RXCDRFREQRESET_IN;
  assign #(in_delay) RXCDRHOLD_INDELAY = RXCDRHOLD_IN;
  assign #(in_delay) RXCDROVRDEN_INDELAY = RXCDROVRDEN_IN;
  assign #(in_delay) RXCDRRESETRSV_INDELAY = RXCDRRESETRSV_IN;
  assign #(in_delay) RXCDRRESET_INDELAY = RXCDRRESET_IN;
  assign #(in_delay) RXCHBONDEN_INDELAY = RXCHBONDEN_IN;
  assign #(in_delay) RXCHBONDI_INDELAY = RXCHBONDI_IN;
  assign #(in_delay) RXCHBONDLEVEL_INDELAY = RXCHBONDLEVEL_IN;
  assign #(in_delay) RXCHBONDMASTER_INDELAY = RXCHBONDMASTER_IN;
  assign #(in_delay) RXCHBONDSLAVE_INDELAY = RXCHBONDSLAVE_IN;
  assign #(in_delay) RXCOMMADETEN_INDELAY = RXCOMMADETEN_IN;
  assign #(in_delay) RXDDIEN_INDELAY = RXDDIEN_IN;
  assign #(in_delay) RXDFEAGCHOLD_INDELAY = RXDFEAGCHOLD_IN;
  assign #(in_delay) RXDFEAGCOVRDEN_INDELAY = RXDFEAGCOVRDEN_IN;
  assign #(in_delay) RXDFECM1EN_INDELAY = RXDFECM1EN_IN;
  assign #(in_delay) RXDFELFHOLD_INDELAY = RXDFELFHOLD_IN;
  assign #(in_delay) RXDFELFOVRDEN_INDELAY = RXDFELFOVRDEN_IN;
  assign #(in_delay) RXDFELPMRESET_INDELAY = RXDFELPMRESET_IN;
  assign #(in_delay) RXDFETAP2HOLD_INDELAY = RXDFETAP2HOLD_IN;
  assign #(in_delay) RXDFETAP2OVRDEN_INDELAY = RXDFETAP2OVRDEN_IN;
  assign #(in_delay) RXDFETAP3HOLD_INDELAY = RXDFETAP3HOLD_IN;
  assign #(in_delay) RXDFETAP3OVRDEN_INDELAY = RXDFETAP3OVRDEN_IN;
  assign #(in_delay) RXDFETAP4HOLD_INDELAY = RXDFETAP4HOLD_IN;
  assign #(in_delay) RXDFETAP4OVRDEN_INDELAY = RXDFETAP4OVRDEN_IN;
  assign #(in_delay) RXDFETAP5HOLD_INDELAY = RXDFETAP5HOLD_IN;
  assign #(in_delay) RXDFETAP5OVRDEN_INDELAY = RXDFETAP5OVRDEN_IN;
  assign #(in_delay) RXDFEUTHOLD_INDELAY = RXDFEUTHOLD_IN;
  assign #(in_delay) RXDFEUTOVRDEN_INDELAY = RXDFEUTOVRDEN_IN;
  assign #(in_delay) RXDFEVPHOLD_INDELAY = RXDFEVPHOLD_IN;
  assign #(in_delay) RXDFEVPOVRDEN_INDELAY = RXDFEVPOVRDEN_IN;
  assign #(in_delay) RXDFEVSEN_INDELAY = RXDFEVSEN_IN;
  assign #(in_delay) RXDFEXYDEN_INDELAY = RXDFEXYDEN_IN;
  assign #(in_delay) RXDFEXYDHOLD_INDELAY = RXDFEXYDHOLD_IN;
  assign #(in_delay) RXDFEXYDOVRDEN_INDELAY = RXDFEXYDOVRDEN_IN;
  assign #(in_delay) RXDLYBYPASS_INDELAY = RXDLYBYPASS_IN;
  assign #(in_delay) RXDLYEN_INDELAY = RXDLYEN_IN;
  assign #(in_delay) RXDLYOVRDEN_INDELAY = RXDLYOVRDEN_IN;
  assign #(in_delay) RXDLYSRESET_INDELAY = RXDLYSRESET_IN;
  assign #(in_delay) RXELECIDLEMODE_INDELAY = RXELECIDLEMODE_IN;
  assign #(in_delay) RXGEARBOXSLIP_INDELAY = RXGEARBOXSLIP_IN;
  assign #(in_delay) RXLPMEN_INDELAY = RXLPMEN_IN;
  assign #(in_delay) RXLPMHFHOLD_INDELAY = RXLPMHFHOLD_IN;
  assign #(in_delay) RXLPMHFOVRDEN_INDELAY = RXLPMHFOVRDEN_IN;
  assign #(in_delay) RXLPMLFHOLD_INDELAY = RXLPMLFHOLD_IN;
  assign #(in_delay) RXLPMLFKLOVRDEN_INDELAY = RXLPMLFKLOVRDEN_IN;
  assign #(in_delay) RXMCOMMAALIGNEN_INDELAY = RXMCOMMAALIGNEN_IN;
  assign #(in_delay) RXMONITORSEL_INDELAY = RXMONITORSEL_IN;
  assign #(in_delay) RXOOBRESET_INDELAY = RXOOBRESET_IN;
  assign #(in_delay) RXOSHOLD_INDELAY = RXOSHOLD_IN;
  assign #(in_delay) RXOSOVRDEN_INDELAY = RXOSOVRDEN_IN;
  assign #(in_delay) RXOUTCLKSEL_INDELAY = RXOUTCLKSEL_IN;
  assign #(in_delay) RXPCOMMAALIGNEN_INDELAY = RXPCOMMAALIGNEN_IN;
  assign #(in_delay) RXPCSRESET_INDELAY = RXPCSRESET_IN;
  assign #(in_delay) RXPD_INDELAY = RXPD_IN;
  assign #(in_delay) RXPHALIGNEN_INDELAY = RXPHALIGNEN_IN;
  assign #(in_delay) RXPHALIGN_INDELAY = RXPHALIGN_IN;
  assign #(in_delay) RXPHDLYPD_INDELAY = RXPHDLYPD_IN;
  assign #(in_delay) RXPHDLYRESET_INDELAY = RXPHDLYRESET_IN;
  assign #(in_delay) RXPHOVRDEN_INDELAY = RXPHOVRDEN_IN;
  assign #(in_delay) RXPMARESET_INDELAY = RXPMARESET_IN;
  assign #(in_delay) RXPOLARITY_INDELAY = RXPOLARITY_IN;
  assign #(in_delay) RXPRBSCNTRESET_INDELAY = RXPRBSCNTRESET_IN;
  assign #(in_delay) RXPRBSSEL_INDELAY = RXPRBSSEL_IN;
  assign #(in_delay) RXQPIEN_INDELAY = RXQPIEN_IN;
  assign #(in_delay) RXRATE_INDELAY = RXRATE_IN;
  assign #(in_delay) RXSLIDE_INDELAY = RXSLIDE_IN;
  assign #(in_delay) RXSYSCLKSEL_INDELAY = RXSYSCLKSEL_IN;
  assign #(in_delay) RXUSERRDY_INDELAY = RXUSERRDY_IN;
  assign #(in_delay) SETERRSTATUS_INDELAY = SETERRSTATUS_IN;
  assign #(in_delay) TSTIN_INDELAY = TSTIN_IN;
  assign #(in_delay) TX8B10BBYPASS_INDELAY = TX8B10BBYPASS_IN;
  assign #(in_delay) TX8B10BEN_INDELAY = TX8B10BEN_IN;
  assign #(in_delay) TXBUFDIFFCTRL_INDELAY = TXBUFDIFFCTRL_IN;
  assign #(in_delay) TXCHARDISPMODE_INDELAY = TXCHARDISPMODE_IN;
  assign #(in_delay) TXCHARDISPVAL_INDELAY = TXCHARDISPVAL_IN;
  assign #(in_delay) TXCHARISK_INDELAY = TXCHARISK_IN;
  assign #(in_delay) TXCOMINIT_INDELAY = TXCOMINIT_IN;
  assign #(in_delay) TXCOMSAS_INDELAY = TXCOMSAS_IN;
  assign #(in_delay) TXCOMWAKE_INDELAY = TXCOMWAKE_IN;
  assign #(in_delay) TXDATA_INDELAY = TXDATA_IN;
  assign #(in_delay) TXDEEMPH_INDELAY = TXDEEMPH_IN;
  assign #(in_delay) TXDETECTRX_INDELAY = TXDETECTRX_IN;
  assign #(in_delay) TXDIFFCTRL_INDELAY = TXDIFFCTRL_IN;
  assign #(in_delay) TXDIFFPD_INDELAY = TXDIFFPD_IN;
  assign #(in_delay) TXDLYBYPASS_INDELAY = TXDLYBYPASS_IN;
  assign #(in_delay) TXDLYEN_INDELAY = TXDLYEN_IN;
  assign #(in_delay) TXDLYHOLD_INDELAY = TXDLYHOLD_IN;
  assign #(in_delay) TXDLYOVRDEN_INDELAY = TXDLYOVRDEN_IN;
  assign #(in_delay) TXDLYSRESET_INDELAY = TXDLYSRESET_IN;
  assign #(in_delay) TXDLYUPDOWN_INDELAY = TXDLYUPDOWN_IN;
  assign #(in_delay) TXELECIDLE_INDELAY = TXELECIDLE_IN;
  assign #(in_delay) TXHEADER_INDELAY = TXHEADER_IN;
  assign #(in_delay) TXINHIBIT_INDELAY = TXINHIBIT_IN;
  assign #(in_delay) TXMAINCURSOR_INDELAY = TXMAINCURSOR_IN;
  assign #(in_delay) TXMARGIN_INDELAY = TXMARGIN_IN;
  assign #(in_delay) TXOUTCLKSEL_INDELAY = TXOUTCLKSEL_IN;
  assign #(in_delay) TXPCSRESET_INDELAY = TXPCSRESET_IN;
  assign #(in_delay) TXPDELECIDLEMODE_INDELAY = TXPDELECIDLEMODE_IN;
  assign #(in_delay) TXPD_INDELAY = TXPD_IN;
  assign #(in_delay) TXPHALIGNEN_INDELAY = TXPHALIGNEN_IN;
  assign #(in_delay) TXPHALIGN_INDELAY = TXPHALIGN_IN;
  assign #(in_delay) TXPHDLYPD_INDELAY = TXPHDLYPD_IN;
  assign #(in_delay) TXPHDLYRESET_INDELAY = TXPHDLYRESET_IN;
  assign #(in_delay) TXPHINIT_INDELAY = TXPHINIT_IN;
  assign #(in_delay) TXPHOVRDEN_INDELAY = TXPHOVRDEN_IN;
  assign #(in_delay) TXPISOPD_INDELAY = TXPISOPD_IN;
  assign #(in_delay) TXPMARESET_INDELAY = TXPMARESET_IN;
  assign #(in_delay) TXPOLARITY_INDELAY = TXPOLARITY_IN;
  assign #(in_delay) TXPOSTCURSORINV_INDELAY = TXPOSTCURSORINV_IN;
  assign #(in_delay) TXPOSTCURSOR_INDELAY = TXPOSTCURSOR_IN;
  assign #(in_delay) TXPRBSFORCEERR_INDELAY = TXPRBSFORCEERR_IN;
  assign #(in_delay) TXPRBSSEL_INDELAY = TXPRBSSEL_IN;
  assign #(in_delay) TXPRECURSORINV_INDELAY = TXPRECURSORINV_IN;
  assign #(in_delay) TXPRECURSOR_INDELAY = TXPRECURSOR_IN;
  assign #(in_delay) TXQPIBIASEN_INDELAY = TXQPIBIASEN_IN;
  assign #(in_delay) TXQPISTRONGPDOWN_INDELAY = TXQPISTRONGPDOWN_IN;
  assign #(in_delay) TXQPIWEAKPUP_INDELAY = TXQPIWEAKPUP_IN;
  assign #(in_delay) TXRATE_INDELAY = TXRATE_IN;
  assign #(in_delay) TXSEQUENCE_INDELAY = TXSEQUENCE_IN;
  assign #(in_delay) TXSTARTSEQ_INDELAY = TXSTARTSEQ_IN;
  assign #(in_delay) TXSWING_INDELAY = TXSWING_IN;
  assign #(in_delay) TXSYSCLKSEL_INDELAY = TXSYSCLKSEL_IN;
  assign #(in_delay) TXUSERRDY_INDELAY = TXUSERRDY_IN;
  assign delay_CFGRESET = CFGRESET_INDELAY;
  assign delay_CLKRSVD = CLKRSVD_INDELAY;
  assign delay_CPLLLOCKDETCLK = CPLLLOCKDETCLK_INDELAY;
  assign delay_CPLLLOCKEN = CPLLLOCKEN_INDELAY;
  assign delay_CPLLPD = CPLLPD_INDELAY;
  assign delay_CPLLREFCLKSEL = CPLLREFCLKSEL_INDELAY;
  assign delay_CPLLRESET = CPLLRESET_INDELAY;
  assign delay_EYESCANMODE = EYESCANMODE_INDELAY;
  assign delay_EYESCANRESET = EYESCANRESET_INDELAY;
  assign delay_EYESCANTRIGGER = EYESCANTRIGGER_INDELAY;
  assign delay_GTGREFCLK = GTGREFCLK_INDELAY;
  assign delay_GTNORTHREFCLK0 = GTNORTHREFCLK0_INDELAY;
  assign delay_GTNORTHREFCLK1 = GTNORTHREFCLK1_INDELAY;
  assign delay_GTREFCLK0 = GTREFCLK0_INDELAY;
  assign delay_GTREFCLK1 = GTREFCLK1_INDELAY;
  assign delay_GTRESETSEL = GTRESETSEL_INDELAY;
  assign delay_GTRSVD = GTRSVD_INDELAY;
  assign delay_GTRXRESET = GTRXRESET_INDELAY;
  assign delay_GTSOUTHREFCLK0 = GTSOUTHREFCLK0_INDELAY;
  assign delay_GTSOUTHREFCLK1 = GTSOUTHREFCLK1_INDELAY;
  assign delay_GTTXRESET = GTTXRESET_INDELAY;
  assign delay_GTXRXN = GTXRXN_INDELAY;
  assign delay_GTXRXP = GTXRXP_INDELAY;
  assign delay_LOOPBACK = LOOPBACK_INDELAY;
  assign delay_PCSRSVDIN = PCSRSVDIN_INDELAY;
  assign delay_PCSRSVDIN2 = PCSRSVDIN2_INDELAY;
  assign delay_PMARSVDIN = PMARSVDIN_INDELAY;
  assign delay_PMARSVDIN2 = PMARSVDIN2_INDELAY;
  assign delay_QPLLCLK = QPLLCLK_INDELAY;
  assign delay_QPLLREFCLK = QPLLREFCLK_INDELAY;
  assign delay_RESETOVRD = RESETOVRD_INDELAY;
  assign delay_RXBUFRESET = RXBUFRESET_INDELAY;
  assign delay_RXCDRFREQRESET = RXCDRFREQRESET_INDELAY;
  assign delay_RXCDRHOLD = RXCDRHOLD_INDELAY;
  assign delay_RXCDROVRDEN = RXCDROVRDEN_INDELAY;
  assign delay_RXCDRRESET = RXCDRRESET_INDELAY;
  assign delay_RXCDRRESETRSV = RXCDRRESETRSV_INDELAY;
  assign delay_RXCHBONDI = RXCHBONDI_INDELAY;
  assign delay_RXDDIEN = RXDDIEN_INDELAY;
  assign delay_RXDFEAGCHOLD = RXDFEAGCHOLD_INDELAY;
  assign delay_RXDFEAGCOVRDEN = RXDFEAGCOVRDEN_INDELAY;
  assign delay_RXDFECM1EN = RXDFECM1EN_INDELAY;
  assign delay_RXDFELFHOLD = RXDFELFHOLD_INDELAY;
  assign delay_RXDFELFOVRDEN = RXDFELFOVRDEN_INDELAY;
  assign delay_RXDFELPMRESET = RXDFELPMRESET_INDELAY;
  assign delay_RXDFETAP2HOLD = RXDFETAP2HOLD_INDELAY;
  assign delay_RXDFETAP2OVRDEN = RXDFETAP2OVRDEN_INDELAY;
  assign delay_RXDFETAP3HOLD = RXDFETAP3HOLD_INDELAY;
  assign delay_RXDFETAP3OVRDEN = RXDFETAP3OVRDEN_INDELAY;
  assign delay_RXDFETAP4HOLD = RXDFETAP4HOLD_INDELAY;
  assign delay_RXDFETAP4OVRDEN = RXDFETAP4OVRDEN_INDELAY;
  assign delay_RXDFETAP5HOLD = RXDFETAP5HOLD_INDELAY;
  assign delay_RXDFETAP5OVRDEN = RXDFETAP5OVRDEN_INDELAY;
  assign delay_RXDFEUTHOLD = RXDFEUTHOLD_INDELAY;
  assign delay_RXDFEUTOVRDEN = RXDFEUTOVRDEN_INDELAY;
  assign delay_RXDFEVPHOLD = RXDFEVPHOLD_INDELAY;
  assign delay_RXDFEVPOVRDEN = RXDFEVPOVRDEN_INDELAY;
  assign delay_RXDFEVSEN = RXDFEVSEN_INDELAY;
  assign delay_RXDFEXYDEN = RXDFEXYDEN_INDELAY;
  assign delay_RXDFEXYDHOLD = RXDFEXYDHOLD_INDELAY;
  assign delay_RXDFEXYDOVRDEN = RXDFEXYDOVRDEN_INDELAY;
  assign delay_RXDLYBYPASS = RXDLYBYPASS_INDELAY;
  assign delay_RXDLYEN = RXDLYEN_INDELAY;
  assign delay_RXDLYOVRDEN = RXDLYOVRDEN_INDELAY;
  assign delay_RXDLYSRESET = RXDLYSRESET_INDELAY;
  assign delay_RXELECIDLEMODE = RXELECIDLEMODE_INDELAY;
  assign delay_RXLPMEN = RXLPMEN_INDELAY;
  assign delay_RXLPMHFHOLD = RXLPMHFHOLD_INDELAY;
  assign delay_RXLPMHFOVRDEN = RXLPMHFOVRDEN_INDELAY;
  assign delay_RXLPMLFHOLD = RXLPMLFHOLD_INDELAY;
  assign delay_RXLPMLFKLOVRDEN = RXLPMLFKLOVRDEN_INDELAY;
  assign delay_RXMONITORSEL = RXMONITORSEL_INDELAY;
  assign delay_RXOOBRESET = RXOOBRESET_INDELAY;
  assign delay_RXOSHOLD = RXOSHOLD_INDELAY;
  assign delay_RXOSOVRDEN = RXOSOVRDEN_INDELAY;
  assign delay_RXOUTCLKSEL = RXOUTCLKSEL_INDELAY;
  assign delay_RXPCSRESET = RXPCSRESET_INDELAY;
  assign delay_RXPHALIGN = RXPHALIGN_INDELAY;
  assign delay_RXPHALIGNEN = RXPHALIGNEN_INDELAY;
  assign delay_RXPHDLYPD = RXPHDLYPD_INDELAY;
  assign delay_RXPHDLYRESET = RXPHDLYRESET_INDELAY;
  assign delay_RXPHOVRDEN = RXPHOVRDEN_INDELAY;
  assign delay_RXPMARESET = RXPMARESET_INDELAY;
  assign delay_RXQPIEN = RXQPIEN_INDELAY;
  assign delay_RXSYSCLKSEL = RXSYSCLKSEL_INDELAY;
  assign delay_RXUSERRDY = RXUSERRDY_INDELAY;
  assign delay_RXUSRCLK = RXUSRCLK_INDELAY;
  assign delay_TSTIN = TSTIN_INDELAY;
  assign delay_TXBUFDIFFCTRL = TXBUFDIFFCTRL_INDELAY;
  assign delay_TXDEEMPH = TXDEEMPH_INDELAY;
  assign delay_TXDIFFCTRL = TXDIFFCTRL_INDELAY;
  assign delay_TXDIFFPD = TXDIFFPD_INDELAY;
  assign delay_TXDLYBYPASS = TXDLYBYPASS_INDELAY;
  assign delay_TXDLYEN = TXDLYEN_INDELAY;
  assign delay_TXDLYOVRDEN = TXDLYOVRDEN_INDELAY;
  assign delay_TXDLYSRESET = TXDLYSRESET_INDELAY;
  assign delay_TXMAINCURSOR = TXMAINCURSOR_INDELAY;
  assign delay_TXOUTCLKSEL = TXOUTCLKSEL_INDELAY;
  assign delay_TXPCSRESET = TXPCSRESET_INDELAY;
  assign delay_TXPDELECIDLEMODE = TXPDELECIDLEMODE_INDELAY;
  assign delay_TXPHALIGN = TXPHALIGN_INDELAY;
  assign delay_TXPHALIGNEN = TXPHALIGNEN_INDELAY;
  assign delay_TXPHDLYPD = TXPHDLYPD_INDELAY;
  assign delay_TXPHDLYRESET = TXPHDLYRESET_INDELAY;
  assign delay_TXPHINIT = TXPHINIT_INDELAY;
  assign delay_TXPHOVRDEN = TXPHOVRDEN_INDELAY;
  assign delay_TXPISOPD = TXPISOPD_INDELAY;
  assign delay_TXPMARESET = TXPMARESET_INDELAY;
  assign delay_TXPOSTCURSOR = TXPOSTCURSOR_INDELAY;
  assign delay_TXPOSTCURSORINV = TXPOSTCURSORINV_INDELAY;
  assign delay_TXPRECURSOR = TXPRECURSOR_INDELAY;
  assign delay_TXPRECURSORINV = TXPRECURSORINV_INDELAY;
  assign delay_TXQPIBIASEN = TXQPIBIASEN_INDELAY;
  assign delay_TXQPISTRONGPDOWN = TXQPISTRONGPDOWN_INDELAY;
  assign delay_TXQPIWEAKPUP = TXQPIWEAKPUP_INDELAY;
  assign delay_TXSYSCLKSEL = TXSYSCLKSEL_INDELAY;
  assign delay_TXUSERRDY = TXUSERRDY_INDELAY;
  assign delay_TXUSRCLK = TXUSRCLK_INDELAY;

  B_GTXE2_CHANNEL #(
    .ALIGN_COMMA_DOUBLE (ALIGN_COMMA_DOUBLE),
    .ALIGN_COMMA_ENABLE (ALIGN_COMMA_ENABLE),
    .ALIGN_COMMA_WORD (ALIGN_COMMA_WORD),
    .ALIGN_MCOMMA_DET (ALIGN_MCOMMA_DET),
    .ALIGN_MCOMMA_VALUE (ALIGN_MCOMMA_VALUE),
    .ALIGN_PCOMMA_DET (ALIGN_PCOMMA_DET),
    .ALIGN_PCOMMA_VALUE (ALIGN_PCOMMA_VALUE),
    .CBCC_DATA_SOURCE_SEL (CBCC_DATA_SOURCE_SEL),
    .CHAN_BOND_KEEP_ALIGN (CHAN_BOND_KEEP_ALIGN),
    .CHAN_BOND_MAX_SKEW (CHAN_BOND_MAX_SKEW),
    .CHAN_BOND_SEQ_1_1 (CHAN_BOND_SEQ_1_1),
    .CHAN_BOND_SEQ_1_2 (CHAN_BOND_SEQ_1_2),
    .CHAN_BOND_SEQ_1_3 (CHAN_BOND_SEQ_1_3),
    .CHAN_BOND_SEQ_1_4 (CHAN_BOND_SEQ_1_4),
    .CHAN_BOND_SEQ_1_ENABLE (CHAN_BOND_SEQ_1_ENABLE),
    .CHAN_BOND_SEQ_2_1 (CHAN_BOND_SEQ_2_1),
    .CHAN_BOND_SEQ_2_2 (CHAN_BOND_SEQ_2_2),
    .CHAN_BOND_SEQ_2_3 (CHAN_BOND_SEQ_2_3),
    .CHAN_BOND_SEQ_2_4 (CHAN_BOND_SEQ_2_4),
    .CHAN_BOND_SEQ_2_ENABLE (CHAN_BOND_SEQ_2_ENABLE),
    .CHAN_BOND_SEQ_2_USE (CHAN_BOND_SEQ_2_USE),
    .CHAN_BOND_SEQ_LEN (CHAN_BOND_SEQ_LEN),
    .CLK_CORRECT_USE (CLK_CORRECT_USE),
    .CLK_COR_KEEP_IDLE (CLK_COR_KEEP_IDLE),
    .CLK_COR_MAX_LAT (CLK_COR_MAX_LAT),
    .CLK_COR_MIN_LAT (CLK_COR_MIN_LAT),
    .CLK_COR_PRECEDENCE (CLK_COR_PRECEDENCE),
    .CLK_COR_REPEAT_WAIT (CLK_COR_REPEAT_WAIT),
    .CLK_COR_SEQ_1_1 (CLK_COR_SEQ_1_1),
    .CLK_COR_SEQ_1_2 (CLK_COR_SEQ_1_2),
    .CLK_COR_SEQ_1_3 (CLK_COR_SEQ_1_3),
    .CLK_COR_SEQ_1_4 (CLK_COR_SEQ_1_4),
    .CLK_COR_SEQ_1_ENABLE (CLK_COR_SEQ_1_ENABLE),
    .CLK_COR_SEQ_2_1 (CLK_COR_SEQ_2_1),
    .CLK_COR_SEQ_2_2 (CLK_COR_SEQ_2_2),
    .CLK_COR_SEQ_2_3 (CLK_COR_SEQ_2_3),
    .CLK_COR_SEQ_2_4 (CLK_COR_SEQ_2_4),
    .CLK_COR_SEQ_2_ENABLE (CLK_COR_SEQ_2_ENABLE),
    .CLK_COR_SEQ_2_USE (CLK_COR_SEQ_2_USE),
    .CLK_COR_SEQ_LEN (CLK_COR_SEQ_LEN),
    .CPLL_CFG (CPLL_CFG),
    .CPLL_FBDIV (CPLL_FBDIV),
    .CPLL_FBDIV_45 (CPLL_FBDIV_45),
    .CPLL_INIT_CFG (CPLL_INIT_CFG),
    .CPLL_LOCK_CFG (CPLL_LOCK_CFG),
    .CPLL_REFCLK_DIV (CPLL_REFCLK_DIV),
    .CPLL_RXOUT_DIV (CPLL_RXOUT_DIV),
    .CPLL_TXOUT_DIV (CPLL_TXOUT_DIV),
    .DEC_MCOMMA_DETECT (DEC_MCOMMA_DETECT),
    .DEC_PCOMMA_DETECT (DEC_PCOMMA_DETECT),
    .DEC_VALID_COMMA_ONLY (DEC_VALID_COMMA_ONLY),
    .DMONITOR_CFG (DMONITOR_CFG),
    .ES_CONTROL (ES_CONTROL),
    .ES_ERRDET_EN (ES_ERRDET_EN),
    .ES_EYE_SCAN_EN (ES_EYE_SCAN_EN),
    .ES_HORZ_OFFSET (ES_HORZ_OFFSET),
    .ES_PMA_CFG (ES_PMA_CFG),
    .ES_PRESCALE (ES_PRESCALE),
    .ES_QUALIFIER (ES_QUALIFIER),
    .ES_QUAL_MASK (ES_QUAL_MASK),
    .ES_SDATA_MASK (ES_SDATA_MASK),
    .ES_VERT_OFFSET (ES_VERT_OFFSET),
    .FTS_DESKEW_SEQ_ENABLE (FTS_DESKEW_SEQ_ENABLE),
    .FTS_LANE_DESKEW_CFG (FTS_LANE_DESKEW_CFG),
    .FTS_LANE_DESKEW_EN (FTS_LANE_DESKEW_EN),
    .GEARBOX_MODE (GEARBOX_MODE),
    .OUTREFCLK_SEL_INV (OUTREFCLK_SEL_INV),
    .PCS_PCIE_EN (PCS_PCIE_EN),
    .PCS_RSVD_ATTR (PCS_RSVD_ATTR),
    .PD_TRANS_TIME_FROM_P2 (PD_TRANS_TIME_FROM_P2),
    .PD_TRANS_TIME_NONE_P2 (PD_TRANS_TIME_NONE_P2),
    .PD_TRANS_TIME_TO_P2 (PD_TRANS_TIME_TO_P2),
    .PMA_RSV (PMA_RSV),
    .PMA_RSV2 (PMA_RSV2),
    .PMA_RSV3 (PMA_RSV3),
    .RXBUFRESET_TIME (RXBUFRESET_TIME),
    .RXBUF_ADDR_MODE (RXBUF_ADDR_MODE),
    .RXBUF_EIDLE_HI_CNT (RXBUF_EIDLE_HI_CNT),
    .RXBUF_EIDLE_LO_CNT (RXBUF_EIDLE_LO_CNT),
    .RXBUF_EN (RXBUF_EN),
    .RXBUF_RESET_ON_CB_CHANGE (RXBUF_RESET_ON_CB_CHANGE),
    .RXBUF_RESET_ON_COMMAALIGN (RXBUF_RESET_ON_COMMAALIGN),
    .RXBUF_RESET_ON_EIDLE (RXBUF_RESET_ON_EIDLE),
    .RXBUF_RESET_ON_RATE_CHANGE (RXBUF_RESET_ON_RATE_CHANGE),
    .RXBUF_THRESH_OVFLW (RXBUF_THRESH_OVFLW),
    .RXBUF_THRESH_OVRD (RXBUF_THRESH_OVRD),
    .RXBUF_THRESH_UNDFLW (RXBUF_THRESH_UNDFLW),
    .RXCDRFREQRESET_TIME (RXCDRFREQRESET_TIME),
    .RXCDRPHRESET_TIME (RXCDRPHRESET_TIME),
    .RXCDR_CFG (RXCDR_CFG),
    .RXCDR_FR_RESET_ON_EIDLE (RXCDR_FR_RESET_ON_EIDLE),
    .RXCDR_HOLD_DURING_EIDLE (RXCDR_HOLD_DURING_EIDLE),
    .RXCDR_LOCK_CFG (RXCDR_LOCK_CFG),
    .RXCDR_PH_RESET_ON_EIDLE (RXCDR_PH_RESET_ON_EIDLE),
    .RXDFELPMRESET_TIME (RXDFELPMRESET_TIME),
    .RXDLY_CFG (RXDLY_CFG),
    .RXDLY_LCFG (RXDLY_LCFG),
    .RXDLY_TAP_CFG (RXDLY_TAP_CFG),
    .RXGEARBOX_EN (RXGEARBOX_EN),
    .RXISCANRESET_TIME (RXISCANRESET_TIME),
    .RXLPM_HF_CFG (RXLPM_HF_CFG),
    .RXLPM_LF_CFG (RXLPM_LF_CFG),
    .RXOOB_CFG (RXOOB_CFG),
    .RXPCSRESET_TIME (RXPCSRESET_TIME),
    .RXPHDLY_CFG (RXPHDLY_CFG),
    .RXPH_CFG (RXPH_CFG),
    .RXPH_MONITOR_SEL (RXPH_MONITOR_SEL),
    .RXPMARESET_TIME (RXPMARESET_TIME),
    .RXPRBS_ERR_LOOPBACK (RXPRBS_ERR_LOOPBACK),
    .RXSLIDE_AUTO_WAIT (RXSLIDE_AUTO_WAIT),
    .RXSLIDE_MODE (RXSLIDE_MODE),
    .RX_BIAS_CFG (RX_BIAS_CFG),
    .RX_BUFFER_CFG (RX_BUFFER_CFG),
    .RX_CLK25_DIV (RX_CLK25_DIV),
    .RX_CLKMUX_PD (RX_CLKMUX_PD),
    .RX_CM_SEL (RX_CM_SEL),
    .RX_CM_TRIM (RX_CM_TRIM),
    .RX_DATA_WIDTH (RX_DATA_WIDTH),
    .RX_DDI_SEL (RX_DDI_SEL),
    .RX_DEBUG_CFG (RX_DEBUG_CFG),
    .RX_DEFER_RESET_BUF_EN (RX_DEFER_RESET_BUF_EN),
    .RX_DFE_GAIN_CFG (RX_DFE_GAIN_CFG),
    .RX_DFE_H2_CFG (RX_DFE_H2_CFG),
    .RX_DFE_H3_CFG (RX_DFE_H3_CFG),
    .RX_DFE_H4_CFG (RX_DFE_H4_CFG),
    .RX_DFE_H5_CFG (RX_DFE_H5_CFG),
    .RX_DFE_KL_CFG (RX_DFE_KL_CFG),
    .RX_DFE_LPM_CFG (RX_DFE_LPM_CFG),
    .RX_DFE_LPM_HOLD_DURING_EIDLE (RX_DFE_LPM_HOLD_DURING_EIDLE),
    .RX_DFE_UT_CFG (RX_DFE_UT_CFG),
    .RX_DFE_VP_CFG (RX_DFE_VP_CFG),
    .RX_DFE_XYD_CFG (RX_DFE_XYD_CFG),
    .RX_DISPERR_SEQ_MATCH (RX_DISPERR_SEQ_MATCH),
    .RX_INT_DATAWIDTH (RX_INT_DATAWIDTH),
    .RX_OS_CFG (RX_OS_CFG),
    .RX_SIG_VALID_DLY (RX_SIG_VALID_DLY),
    .RX_XCLK_SEL (RX_XCLK_SEL),
    .SAS_MAX_COM (SAS_MAX_COM),
    .SAS_MIN_COM (SAS_MIN_COM),
    .SATA_BURST_SEQ_LEN (SATA_BURST_SEQ_LEN),
    .SATA_BURST_VAL (SATA_BURST_VAL),
    .SATA_CPLL_CFG (SATA_CPLL_CFG),
    .SATA_EIDLE_VAL (SATA_EIDLE_VAL),
    .SATA_MAX_BURST (SATA_MAX_BURST),
    .SATA_MAX_INIT (SATA_MAX_INIT),
    .SATA_MAX_WAKE (SATA_MAX_WAKE),
    .SATA_MIN_BURST (SATA_MIN_BURST),
    .SATA_MIN_INIT (SATA_MIN_INIT),
    .SATA_MIN_WAKE (SATA_MIN_WAKE),
    .SHOW_REALIGN_COMMA (SHOW_REALIGN_COMMA),
    .SIM_CPLLREFCLK_SEL (SIM_CPLLREFCLK_SEL),
    .SIM_RECEIVER_DETECT_PASS (SIM_RECEIVER_DETECT_PASS),
    .SIM_RESET_SPEEDUP (SIM_RESET_SPEEDUP),
    .SIM_TX_EIDLE_DRIVE_LEVEL (SIM_TX_EIDLE_DRIVE_LEVEL),
    .SIM_VERSION (SIM_VERSION),
    .TERM_RCAL_CFG (TERM_RCAL_CFG),
    .TERM_RCAL_OVRD (TERM_RCAL_OVRD),
    .TRANS_TIME_RATE (TRANS_TIME_RATE),
    .TST_RSV (TST_RSV),
    .TXBUF_EN (TXBUF_EN),
    .TXBUF_RESET_ON_RATE_CHANGE (TXBUF_RESET_ON_RATE_CHANGE),
    .TXDLY_CFG (TXDLY_CFG),
    .TXDLY_LCFG (TXDLY_LCFG),
    .TXDLY_TAP_CFG (TXDLY_TAP_CFG),
    .TXGEARBOX_EN (TXGEARBOX_EN),
    .TXPCSRESET_TIME (TXPCSRESET_TIME),
    .TXPHDLY_CFG (TXPHDLY_CFG),
    .TXPH_CFG (TXPH_CFG),
    .TXPH_MONITOR_SEL (TXPH_MONITOR_SEL),
    .TXPMARESET_TIME (TXPMARESET_TIME),
    .TX_CLK25_DIV (TX_CLK25_DIV),
    .TX_CLKMUX_PD (TX_CLKMUX_PD),
    .TX_DATA_WIDTH (TX_DATA_WIDTH),
    .TX_DEEMPH0 (TX_DEEMPH0),
    .TX_DEEMPH1 (TX_DEEMPH1),
    .TX_DRIVE_MODE (TX_DRIVE_MODE),
    .TX_EIDLE_ASSERT_DELAY (TX_EIDLE_ASSERT_DELAY),
    .TX_EIDLE_DEASSERT_DELAY (TX_EIDLE_DEASSERT_DELAY),
    .TX_INT_DATAWIDTH (TX_INT_DATAWIDTH),
    .TX_LOOPBACK_DRIVE_HIZ (TX_LOOPBACK_DRIVE_HIZ),
    .TX_MAINCURSOR_SEL (TX_MAINCURSOR_SEL),
    .TX_MARGIN_FULL_0 (TX_MARGIN_FULL_0),
    .TX_MARGIN_FULL_1 (TX_MARGIN_FULL_1),
    .TX_MARGIN_FULL_2 (TX_MARGIN_FULL_2),
    .TX_MARGIN_FULL_3 (TX_MARGIN_FULL_3),
    .TX_MARGIN_FULL_4 (TX_MARGIN_FULL_4),
    .TX_MARGIN_LOW_0 (TX_MARGIN_LOW_0),
    .TX_MARGIN_LOW_1 (TX_MARGIN_LOW_1),
    .TX_MARGIN_LOW_2 (TX_MARGIN_LOW_2),
    .TX_MARGIN_LOW_3 (TX_MARGIN_LOW_3),
    .TX_MARGIN_LOW_4 (TX_MARGIN_LOW_4),
    .TX_PREDRIVER_MODE (TX_PREDRIVER_MODE),
    .TX_QPI_STATUS_EN (TX_QPI_STATUS_EN),
    .TX_RXDETECT_CFG (TX_RXDETECT_CFG),
    .TX_RXDETECT_REF (TX_RXDETECT_REF),
    .TX_XCLK_SEL (TX_XCLK_SEL),
    .UCODEER_CLR (UCODEER_CLR))

    B_GTXE2_CHANNEL_INST (
    .CPLLFBCLKLOST (delay_CPLLFBCLKLOST),
    .CPLLLOCK (delay_CPLLLOCK),
    .CPLLREFCLKLOST (delay_CPLLREFCLKLOST),
    .DMONITOROUT (delay_DMONITOROUT),
    .DRPDO (delay_DRPDO),
    .DRPRDY (delay_DRPRDY),
    .EYESCANDATAERROR (delay_EYESCANDATAERROR),
    .GTREFCLKMONITOR (delay_GTREFCLKMONITOR),
    .GTXTXN (delay_GTXTXN),
    .GTXTXP (delay_GTXTXP),
    .PCSRSVDOUT (delay_PCSRSVDOUT),
    .PHYSTATUS (delay_PHYSTATUS),
    .RXBUFSTATUS (delay_RXBUFSTATUS),
    .RXBYTEISALIGNED (delay_RXBYTEISALIGNED),
    .RXBYTEREALIGN (delay_RXBYTEREALIGN),
    .RXCDRLOCK (delay_RXCDRLOCK),
    .RXCHANBONDSEQ (delay_RXCHANBONDSEQ),
    .RXCHANISALIGNED (delay_RXCHANISALIGNED),
    .RXCHANREALIGN (delay_RXCHANREALIGN),
    .RXCHARISCOMMA (delay_RXCHARISCOMMA),
    .RXCHARISK (delay_RXCHARISK),
    .RXCHBONDO (delay_RXCHBONDO),
    .RXCLKCORCNT (delay_RXCLKCORCNT),
    .RXCOMINITDET (delay_RXCOMINITDET),
    .RXCOMMADET (delay_RXCOMMADET),
    .RXCOMSASDET (delay_RXCOMSASDET),
    .RXCOMWAKEDET (delay_RXCOMWAKEDET),
    .RXDATA (delay_RXDATA),
    .RXDATAVALID (delay_RXDATAVALID),
    .RXDISPERR (delay_RXDISPERR),
    .RXDLYSRESETDONE (delay_RXDLYSRESETDONE),
    .RXELECIDLE (delay_RXELECIDLE),
    .RXHEADER (delay_RXHEADER),
    .RXHEADERVALID (delay_RXHEADERVALID),
    .RXMONITOROUT (delay_RXMONITOROUT),
    .RXNOTINTABLE (delay_RXNOTINTABLE),
    .RXOUTCLK (delay_RXOUTCLK),
    .RXOUTCLKFABRIC (delay_RXOUTCLKFABRIC),
    .RXOUTCLKPCS (delay_RXOUTCLKPCS),
    .RXPHALIGNDONE (delay_RXPHALIGNDONE),
    .RXPHMONITOR (delay_RXPHMONITOR),
    .RXPHSLIPMONITOR (delay_RXPHSLIPMONITOR),
    .RXPRBSERR (delay_RXPRBSERR),
    .RXQPISENN (delay_RXQPISENN),
    .RXQPISENP (delay_RXQPISENP),
    .RXRATEDONE (delay_RXRATEDONE),
    .RXRESETDONE (delay_RXRESETDONE),
    .RXSTARTOFSEQ (delay_RXSTARTOFSEQ),
    .RXSTATUS (delay_RXSTATUS),
    .RXVALID (delay_RXVALID),
    .TSTOUT (delay_TSTOUT),
    .TXBUFSTATUS (delay_TXBUFSTATUS),
    .TXCOMFINISH (delay_TXCOMFINISH),
    .TXDLYSRESETDONE (delay_TXDLYSRESETDONE),
    .TXGEARBOXREADY (delay_TXGEARBOXREADY),
    .TXOUTCLK (delay_TXOUTCLK),
    .TXOUTCLKFABRIC (delay_TXOUTCLKFABRIC),
    .TXOUTCLKPCS (delay_TXOUTCLKPCS),
    .TXPHALIGNDONE (delay_TXPHALIGNDONE),
    .TXPHINITDONE (delay_TXPHINITDONE),
    .TXQPISENN (delay_TXQPISENN),
    .TXQPISENP (delay_TXQPISENP),
    .TXRATEDONE (delay_TXRATEDONE),
    .TXRESETDONE (delay_TXRESETDONE),
    .CFGRESET (delay_CFGRESET),
    .CLKRSVD (delay_CLKRSVD),
    .CPLLLOCKDETCLK (delay_CPLLLOCKDETCLK),
    .CPLLLOCKEN (delay_CPLLLOCKEN),
    .CPLLPD (delay_CPLLPD),
    .CPLLREFCLKSEL (delay_CPLLREFCLKSEL),
    .CPLLRESET (delay_CPLLRESET),
    .DRPADDR (delay_DRPADDR),
    .DRPCLK (delay_DRPCLK),
    .DRPDI (delay_DRPDI),
    .DRPEN (delay_DRPEN),
    .DRPWE (delay_DRPWE),
    .EYESCANMODE (delay_EYESCANMODE),
    .EYESCANRESET (delay_EYESCANRESET),
    .EYESCANTRIGGER (delay_EYESCANTRIGGER),
    .GTGREFCLK (delay_GTGREFCLK),
    .GTNORTHREFCLK0 (delay_GTNORTHREFCLK0),
    .GTNORTHREFCLK1 (delay_GTNORTHREFCLK1),
    .GTREFCLK0 (delay_GTREFCLK0),
    .GTREFCLK1 (delay_GTREFCLK1),
    .GTRESETSEL (delay_GTRESETSEL),
    .GTRSVD (delay_GTRSVD),
    .GTRXRESET (delay_GTRXRESET),
    .GTSOUTHREFCLK0 (delay_GTSOUTHREFCLK0),
    .GTSOUTHREFCLK1 (delay_GTSOUTHREFCLK1),
    .GTTXRESET (delay_GTTXRESET),
    .GTXRXN (delay_GTXRXN),
    .GTXRXP (delay_GTXRXP),
    .LOOPBACK (delay_LOOPBACK),
    .PCSRSVDIN (delay_PCSRSVDIN),
    .PCSRSVDIN2 (delay_PCSRSVDIN2),
    .PMARSVDIN (delay_PMARSVDIN),
    .PMARSVDIN2 (delay_PMARSVDIN2),
    .QPLLCLK (delay_QPLLCLK),
    .QPLLREFCLK (delay_QPLLREFCLK),
    .RESETOVRD (delay_RESETOVRD),
    .RX8B10BEN (delay_RX8B10BEN),
    .RXBUFRESET (delay_RXBUFRESET),
    .RXCDRFREQRESET (delay_RXCDRFREQRESET),
    .RXCDRHOLD (delay_RXCDRHOLD),
    .RXCDROVRDEN (delay_RXCDROVRDEN),
    .RXCDRRESET (delay_RXCDRRESET),
    .RXCDRRESETRSV (delay_RXCDRRESETRSV),
    .RXCHBONDEN (delay_RXCHBONDEN),
    .RXCHBONDI (delay_RXCHBONDI),
    .RXCHBONDLEVEL (delay_RXCHBONDLEVEL),
    .RXCHBONDMASTER (delay_RXCHBONDMASTER),
    .RXCHBONDSLAVE (delay_RXCHBONDSLAVE),
    .RXCOMMADETEN (delay_RXCOMMADETEN),
    .RXDDIEN (delay_RXDDIEN),
    .RXDFEAGCHOLD (delay_RXDFEAGCHOLD),
    .RXDFEAGCOVRDEN (delay_RXDFEAGCOVRDEN),
    .RXDFECM1EN (delay_RXDFECM1EN),
    .RXDFELFHOLD (delay_RXDFELFHOLD),
    .RXDFELFOVRDEN (delay_RXDFELFOVRDEN),
    .RXDFELPMRESET (delay_RXDFELPMRESET),
    .RXDFETAP2HOLD (delay_RXDFETAP2HOLD),
    .RXDFETAP2OVRDEN (delay_RXDFETAP2OVRDEN),
    .RXDFETAP3HOLD (delay_RXDFETAP3HOLD),
    .RXDFETAP3OVRDEN (delay_RXDFETAP3OVRDEN),
    .RXDFETAP4HOLD (delay_RXDFETAP4HOLD),
    .RXDFETAP4OVRDEN (delay_RXDFETAP4OVRDEN),
    .RXDFETAP5HOLD (delay_RXDFETAP5HOLD),
    .RXDFETAP5OVRDEN (delay_RXDFETAP5OVRDEN),
    .RXDFEUTHOLD (delay_RXDFEUTHOLD),
    .RXDFEUTOVRDEN (delay_RXDFEUTOVRDEN),
    .RXDFEVPHOLD (delay_RXDFEVPHOLD),
    .RXDFEVPOVRDEN (delay_RXDFEVPOVRDEN),
    .RXDFEVSEN (delay_RXDFEVSEN),
    .RXDFEXYDEN (delay_RXDFEXYDEN),
    .RXDFEXYDHOLD (delay_RXDFEXYDHOLD),
    .RXDFEXYDOVRDEN (delay_RXDFEXYDOVRDEN),
    .RXDLYBYPASS (delay_RXDLYBYPASS),
    .RXDLYEN (delay_RXDLYEN),
    .RXDLYOVRDEN (delay_RXDLYOVRDEN),
    .RXDLYSRESET (delay_RXDLYSRESET),
    .RXELECIDLEMODE (delay_RXELECIDLEMODE),
    .RXGEARBOXSLIP (delay_RXGEARBOXSLIP),
    .RXLPMEN (delay_RXLPMEN),
    .RXLPMHFHOLD (delay_RXLPMHFHOLD),
    .RXLPMHFOVRDEN (delay_RXLPMHFOVRDEN),
    .RXLPMLFHOLD (delay_RXLPMLFHOLD),
    .RXLPMLFKLOVRDEN (delay_RXLPMLFKLOVRDEN),
    .RXMCOMMAALIGNEN (delay_RXMCOMMAALIGNEN),
    .RXMONITORSEL (delay_RXMONITORSEL),
    .RXOOBRESET (delay_RXOOBRESET),
    .RXOSHOLD (delay_RXOSHOLD),
    .RXOSOVRDEN (delay_RXOSOVRDEN),
    .RXOUTCLKSEL (delay_RXOUTCLKSEL),
    .RXPCOMMAALIGNEN (delay_RXPCOMMAALIGNEN),
    .RXPCSRESET (delay_RXPCSRESET),
    .RXPD (delay_RXPD),
    .RXPHALIGN (delay_RXPHALIGN),
    .RXPHALIGNEN (delay_RXPHALIGNEN),
    .RXPHDLYPD (delay_RXPHDLYPD),
    .RXPHDLYRESET (delay_RXPHDLYRESET),
    .RXPHOVRDEN (delay_RXPHOVRDEN),
    .RXPMARESET (delay_RXPMARESET),
    .RXPOLARITY (delay_RXPOLARITY),
    .RXPRBSCNTRESET (delay_RXPRBSCNTRESET),
    .RXPRBSSEL (delay_RXPRBSSEL),
    .RXQPIEN (delay_RXQPIEN),
    .RXRATE (delay_RXRATE),
    .RXSLIDE (delay_RXSLIDE),
    .RXSYSCLKSEL (delay_RXSYSCLKSEL),
    .RXUSERRDY (delay_RXUSERRDY),
    .RXUSRCLK (delay_RXUSRCLK),
    .RXUSRCLK2 (delay_RXUSRCLK2),
    .SETERRSTATUS (delay_SETERRSTATUS),
    .TSTIN (delay_TSTIN),
    .TX8B10BBYPASS (delay_TX8B10BBYPASS),
    .TX8B10BEN (delay_TX8B10BEN),
    .TXBUFDIFFCTRL (delay_TXBUFDIFFCTRL),
    .TXCHARDISPMODE (delay_TXCHARDISPMODE),
    .TXCHARDISPVAL (delay_TXCHARDISPVAL),
    .TXCHARISK (delay_TXCHARISK),
    .TXCOMINIT (delay_TXCOMINIT),
    .TXCOMSAS (delay_TXCOMSAS),
    .TXCOMWAKE (delay_TXCOMWAKE),
    .TXDATA (delay_TXDATA),
    .TXDEEMPH (delay_TXDEEMPH),
    .TXDETECTRX (delay_TXDETECTRX),
    .TXDIFFCTRL (delay_TXDIFFCTRL),
    .TXDIFFPD (delay_TXDIFFPD),
    .TXDLYBYPASS (delay_TXDLYBYPASS),
    .TXDLYEN (delay_TXDLYEN),
    .TXDLYHOLD (delay_TXDLYHOLD),
    .TXDLYOVRDEN (delay_TXDLYOVRDEN),
    .TXDLYSRESET (delay_TXDLYSRESET),
    .TXDLYUPDOWN (delay_TXDLYUPDOWN),
    .TXELECIDLE (delay_TXELECIDLE),
    .TXHEADER (delay_TXHEADER),
    .TXINHIBIT (delay_TXINHIBIT),
    .TXMAINCURSOR (delay_TXMAINCURSOR),
    .TXMARGIN (delay_TXMARGIN),
    .TXOUTCLKSEL (delay_TXOUTCLKSEL),
    .TXPCSRESET (delay_TXPCSRESET),
    .TXPD (delay_TXPD),
    .TXPDELECIDLEMODE (delay_TXPDELECIDLEMODE),
    .TXPHALIGN (delay_TXPHALIGN),
    .TXPHALIGNEN (delay_TXPHALIGNEN),
    .TXPHDLYPD (delay_TXPHDLYPD),
    .TXPHDLYRESET (delay_TXPHDLYRESET),
    .TXPHDLYTSTCLK (delay_TXPHDLYTSTCLK),
    .TXPHINIT (delay_TXPHINIT),
    .TXPHOVRDEN (delay_TXPHOVRDEN),
    .TXPISOPD (delay_TXPISOPD),
    .TXPMARESET (delay_TXPMARESET),
    .TXPOLARITY (delay_TXPOLARITY),
    .TXPOSTCURSOR (delay_TXPOSTCURSOR),
    .TXPOSTCURSORINV (delay_TXPOSTCURSORINV),
    .TXPRBSFORCEERR (delay_TXPRBSFORCEERR),
    .TXPRBSSEL (delay_TXPRBSSEL),
    .TXPRECURSOR (delay_TXPRECURSOR),
    .TXPRECURSORINV (delay_TXPRECURSORINV),
    .TXQPIBIASEN (delay_TXQPIBIASEN),
    .TXQPISTRONGPDOWN (delay_TXQPISTRONGPDOWN),
    .TXQPIWEAKPUP (delay_TXQPIWEAKPUP),
    .TXRATE (delay_TXRATE),
    .TXSEQUENCE (delay_TXSEQUENCE),
    .TXSTARTSEQ (delay_TXSTARTSEQ),
    .TXSWING (delay_TXSWING),
    .TXSYSCLKSEL (delay_TXSYSCLKSEL),
    .TXUSERRDY (delay_TXUSERRDY),
    .TXUSRCLK (delay_TXUSRCLK),
    .TXUSRCLK2 (delay_TXUSRCLK2),
    .GSR (GSR)
  );

  specify
    $period (posedge CPLLLOCKDETCLK, 0:0:0, notifier);
    $period (posedge DRPCLK, 0:0:0, notifier);
    $period (posedge GTGREFCLK, 0:0:0, notifier);
    $period (posedge GTNORTHREFCLK0, 0:0:0, notifier);
    $period (posedge GTNORTHREFCLK1, 0:0:0, notifier);
    $period (posedge GTREFCLK0, 0:0:0, notifier);
    $period (posedge GTREFCLK1, 0:0:0, notifier);
    $period (posedge GTREFCLKMONITOR, 0:0:0, notifier);
    $period (posedge GTSOUTHREFCLK0, 0:0:0, notifier);
    $period (posedge GTSOUTHREFCLK1, 0:0:0, notifier);
    $period (posedge QPLLCLK, 0:0:0, notifier);
    $period (posedge RXOUTCLK, 0:0:0, notifier);
    $period (posedge RXOUTCLKFABRIC, 0:0:0, notifier);
    $period (posedge RXOUTCLKPCS, 0:0:0, notifier);
    $period (posedge RXUSRCLK, 0:0:0, notifier);
    $period (posedge RXUSRCLK2, 0:0:0, notifier);
    $period (posedge TXOUTCLK, 0:0:0, notifier);
    $period (posedge TXOUTCLKFABRIC, 0:0:0, notifier);
    $period (posedge TXOUTCLKPCS, 0:0:0, notifier);
    $period (posedge TXPHDLYTSTCLK, 0:0:0, notifier);
    $period (posedge TXUSRCLK, 0:0:0, notifier);
    $period (posedge TXUSRCLK2, 0:0:0, notifier);
    $setuphold (posedge DRPCLK, negedge DRPADDR, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR);
    $setuphold (posedge DRPCLK, negedge DRPDI, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI);
    $setuphold (posedge DRPCLK, negedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, negedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge DRPCLK, posedge DRPADDR, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR);
    $setuphold (posedge DRPCLK, posedge DRPDI, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI);
    $setuphold (posedge DRPCLK, posedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, posedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge RXUSRCLK2, negedge RX8B10BEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RX8B10BEN);
    $setuphold (posedge RXUSRCLK2, negedge RXCHBONDEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDEN);
    $setuphold (posedge RXUSRCLK2, negedge RXCHBONDLEVEL, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDLEVEL);
    $setuphold (posedge RXUSRCLK2, negedge RXCHBONDMASTER, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDMASTER);
    $setuphold (posedge RXUSRCLK2, negedge RXCHBONDSLAVE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDSLAVE);
    $setuphold (posedge RXUSRCLK2, negedge RXCOMMADETEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCOMMADETEN);
    $setuphold (posedge RXUSRCLK2, negedge RXGEARBOXSLIP, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXGEARBOXSLIP);
    $setuphold (posedge RXUSRCLK2, negedge RXMCOMMAALIGNEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXMCOMMAALIGNEN);
    $setuphold (posedge RXUSRCLK2, negedge RXPCOMMAALIGNEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPCOMMAALIGNEN);
    $setuphold (posedge RXUSRCLK2, negedge RXPD, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPD);
    $setuphold (posedge RXUSRCLK2, negedge RXPOLARITY, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPOLARITY);
    $setuphold (posedge RXUSRCLK2, negedge RXPRBSCNTRESET, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPRBSCNTRESET);
    $setuphold (posedge RXUSRCLK2, negedge RXPRBSSEL, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPRBSSEL);
    $setuphold (posedge RXUSRCLK2, negedge RXRATE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXRATE);
    $setuphold (posedge RXUSRCLK2, negedge RXSLIDE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXSLIDE);
    $setuphold (posedge RXUSRCLK2, negedge SETERRSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_SETERRSTATUS);
    $setuphold (posedge RXUSRCLK2, posedge RX8B10BEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RX8B10BEN);
    $setuphold (posedge RXUSRCLK2, posedge RXCHBONDEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDEN);
    $setuphold (posedge RXUSRCLK2, posedge RXCHBONDLEVEL, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDLEVEL);
    $setuphold (posedge RXUSRCLK2, posedge RXCHBONDMASTER, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDMASTER);
    $setuphold (posedge RXUSRCLK2, posedge RXCHBONDSLAVE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCHBONDSLAVE);
    $setuphold (posedge RXUSRCLK2, posedge RXCOMMADETEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXCOMMADETEN);
    $setuphold (posedge RXUSRCLK2, posedge RXGEARBOXSLIP, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXGEARBOXSLIP);
    $setuphold (posedge RXUSRCLK2, posedge RXMCOMMAALIGNEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXMCOMMAALIGNEN);
    $setuphold (posedge RXUSRCLK2, posedge RXPCOMMAALIGNEN, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPCOMMAALIGNEN);
    $setuphold (posedge RXUSRCLK2, posedge RXPD, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPD);
    $setuphold (posedge RXUSRCLK2, posedge RXPOLARITY, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPOLARITY);
    $setuphold (posedge RXUSRCLK2, posedge RXPRBSCNTRESET, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPRBSCNTRESET);
    $setuphold (posedge RXUSRCLK2, posedge RXPRBSSEL, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXPRBSSEL);
    $setuphold (posedge RXUSRCLK2, posedge RXRATE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXRATE);
    $setuphold (posedge RXUSRCLK2, posedge RXSLIDE, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_RXSLIDE);
    $setuphold (posedge RXUSRCLK2, posedge SETERRSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RXUSRCLK2, delay_SETERRSTATUS);
    $setuphold (posedge TXPHDLYTSTCLK, negedge TXDLYHOLD, 0:0:0, 0:0:0, notifier,,, delay_TXPHDLYTSTCLK, delay_TXDLYHOLD);
    $setuphold (posedge TXPHDLYTSTCLK, negedge TXDLYUPDOWN, 0:0:0, 0:0:0, notifier,,, delay_TXPHDLYTSTCLK, delay_TXDLYUPDOWN);
    $setuphold (posedge TXPHDLYTSTCLK, posedge TXDLYHOLD, 0:0:0, 0:0:0, notifier,,, delay_TXPHDLYTSTCLK, delay_TXDLYHOLD);
    $setuphold (posedge TXPHDLYTSTCLK, posedge TXDLYUPDOWN, 0:0:0, 0:0:0, notifier,,, delay_TXPHDLYTSTCLK, delay_TXDLYUPDOWN);
    $setuphold (posedge TXUSRCLK2, negedge TX8B10BBYPASS, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TX8B10BBYPASS);
    $setuphold (posedge TXUSRCLK2, negedge TX8B10BEN, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TX8B10BEN);
    $setuphold (posedge TXUSRCLK2, negedge TXCHARDISPMODE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARDISPMODE);
    $setuphold (posedge TXUSRCLK2, negedge TXCHARDISPVAL, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARDISPVAL);
    $setuphold (posedge TXUSRCLK2, negedge TXCHARISK, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARISK);
    $setuphold (posedge TXUSRCLK2, negedge TXCOMINIT, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMINIT);
    $setuphold (posedge TXUSRCLK2, negedge TXCOMSAS, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMSAS);
    $setuphold (posedge TXUSRCLK2, negedge TXCOMWAKE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMWAKE);
    $setuphold (posedge TXUSRCLK2, negedge TXDATA, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXDATA);
    $setuphold (posedge TXUSRCLK2, negedge TXDETECTRX, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXDETECTRX);
    $setuphold (posedge TXUSRCLK2, negedge TXELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXELECIDLE);
    $setuphold (posedge TXUSRCLK2, negedge TXHEADER, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXHEADER);
    $setuphold (posedge TXUSRCLK2, negedge TXINHIBIT, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXINHIBIT);
    $setuphold (posedge TXUSRCLK2, negedge TXMARGIN, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXMARGIN);
    $setuphold (posedge TXUSRCLK2, negedge TXPD, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPD);
    $setuphold (posedge TXUSRCLK2, negedge TXPOLARITY, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPOLARITY);
    $setuphold (posedge TXUSRCLK2, negedge TXPRBSFORCEERR, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPRBSFORCEERR);
    $setuphold (posedge TXUSRCLK2, negedge TXPRBSSEL, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPRBSSEL);
    $setuphold (posedge TXUSRCLK2, negedge TXRATE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXRATE);
    $setuphold (posedge TXUSRCLK2, negedge TXSEQUENCE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSEQUENCE);
    $setuphold (posedge TXUSRCLK2, negedge TXSTARTSEQ, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSTARTSEQ);
    $setuphold (posedge TXUSRCLK2, negedge TXSWING, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSWING);
    $setuphold (posedge TXUSRCLK2, posedge TX8B10BBYPASS, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TX8B10BBYPASS);
    $setuphold (posedge TXUSRCLK2, posedge TX8B10BEN, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TX8B10BEN);
    $setuphold (posedge TXUSRCLK2, posedge TXCHARDISPMODE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARDISPMODE);
    $setuphold (posedge TXUSRCLK2, posedge TXCHARDISPVAL, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARDISPVAL);
    $setuphold (posedge TXUSRCLK2, posedge TXCHARISK, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCHARISK);
    $setuphold (posedge TXUSRCLK2, posedge TXCOMINIT, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMINIT);
    $setuphold (posedge TXUSRCLK2, posedge TXCOMSAS, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMSAS);
    $setuphold (posedge TXUSRCLK2, posedge TXCOMWAKE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXCOMWAKE);
    $setuphold (posedge TXUSRCLK2, posedge TXDATA, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXDATA);
    $setuphold (posedge TXUSRCLK2, posedge TXDETECTRX, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXDETECTRX);
    $setuphold (posedge TXUSRCLK2, posedge TXELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXELECIDLE);
    $setuphold (posedge TXUSRCLK2, posedge TXHEADER, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXHEADER);
    $setuphold (posedge TXUSRCLK2, posedge TXINHIBIT, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXINHIBIT);
    $setuphold (posedge TXUSRCLK2, posedge TXMARGIN, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXMARGIN);
    $setuphold (posedge TXUSRCLK2, posedge TXPD, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPD);
    $setuphold (posedge TXUSRCLK2, posedge TXPOLARITY, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPOLARITY);
    $setuphold (posedge TXUSRCLK2, posedge TXPRBSFORCEERR, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPRBSFORCEERR);
    $setuphold (posedge TXUSRCLK2, posedge TXPRBSSEL, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXPRBSSEL);
    $setuphold (posedge TXUSRCLK2, posedge TXRATE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXRATE);
    $setuphold (posedge TXUSRCLK2, posedge TXSEQUENCE, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSEQUENCE);
    $setuphold (posedge TXUSRCLK2, posedge TXSTARTSEQ, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSTARTSEQ);
    $setuphold (posedge TXUSRCLK2, posedge TXSWING, 0:0:0, 0:0:0, notifier,,, delay_TXUSRCLK2, delay_TXSWING);
    ( DRPCLK *> DRPDO) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPRDY) = (100:100:100, 100:100:100);
    ( GTNORTHREFCLK0 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( GTNORTHREFCLK1 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( GTREFCLK0 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( GTREFCLK1 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( GTSOUTHREFCLK0 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( GTSOUTHREFCLK1 *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( QPLLCLK *> GTREFCLKMONITOR) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> PHYSTATUS) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXBUFSTATUS) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXBYTEISALIGNED) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXBYTEREALIGN) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHANBONDSEQ) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHANISALIGNED) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHANREALIGN) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHARISCOMMA) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHARISK) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCHBONDO) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCLKCORCNT) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCOMINITDET) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCOMMADET) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCOMSASDET) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXCOMWAKEDET) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXDATA) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXDATAVALID) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXDISPERR) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXHEADER) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXHEADERVALID) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXNOTINTABLE) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXPRBSERR) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXRATEDONE) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXRESETDONE) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXSTARTOFSEQ) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXSTATUS) = (100:100:100, 100:100:100);
    ( RXUSRCLK2 *> RXVALID) = (100:100:100, 100:100:100);
    ( TXUSRCLK2 *> TXBUFSTATUS) = (100:100:100, 100:100:100);
    ( TXUSRCLK2 *> TXCOMFINISH) = (100:100:100, 100:100:100);
    ( TXUSRCLK2 *> TXGEARBOXREADY) = (100:100:100, 100:100:100);
    ( TXUSRCLK2 *> TXRATEDONE) = (100:100:100, 100:100:100);
    ( TXUSRCLK2 *> TXRESETDONE) = (100:100:100, 100:100:100);

    specparam PATHPULSE$ = 0;
  endspecify
endmodule
